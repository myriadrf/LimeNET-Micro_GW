-- factory.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity factory is
	port (
		bridge_0_address     : in    std_logic_vector(20 downto 0) := (others => '0'); -- bridge_0.address
		bridge_0_byte_enable : in    std_logic_vector(3 downto 0)  := (others => '0'); --         .byte_enable
		bridge_0_read        : in    std_logic                     := '0';             --         .read
		bridge_0_write       : in    std_logic                     := '0';             --         .write
		bridge_0_write_data  : in    std_logic_vector(31 downto 0) := (others => '0'); --         .write_data
		bridge_0_acknowledge : out   std_logic;                                        --         .acknowledge
		bridge_0_read_data   : out   std_logic_vector(31 downto 0);                    --         .read_data
		clk_clk              : in    std_logic                     := '0';             --      clk.clk
		extfifo_of_d         : out   std_logic_vector(31 downto 0);                    --  extfifo.of_d
		extfifo_of_wr        : out   std_logic;                                        --         .of_wr
		extfifo_of_wrfull    : in    std_logic                     := '0';             --         .of_wrfull
		extfifo_if_d         : in    std_logic_vector(31 downto 0) := (others => '0'); --         .if_d
		extfifo_if_rd        : out   std_logic;                                        --         .if_rd
		extfifo_if_rdempty   : in    std_logic                     := '0';             --         .if_rdempty
		extfifo_fifo_rst     : out   std_logic;                                        --         .fifo_rst
		pio_0_export         : out   std_logic_vector(7 downto 0);                     --    pio_0.export
		reset_reset_n        : in    std_logic                     := '0';             --    reset.reset_n
		scl_export           : inout std_logic                     := '0';             --      scl.export
		sda_export           : inout std_logic                     := '0'              --      sda.export
	);
end entity factory;

architecture rtl of factory is
	component avs_fifo_int is
		port (
			avs_s0_address     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avs_s0_read        : in  std_logic                     := 'X';             -- read
			avs_s0_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s0_write       : in  std_logic                     := 'X';             -- write
			avs_s0_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s0_waitrequest : out std_logic;                                        -- waitrequest
			clock_clk          : in  std_logic                     := 'X';             -- clk
			reset_reset        : in  std_logic                     := 'X';             -- reset
			of_d               : out std_logic_vector(31 downto 0);                    -- of_d
			of_wr              : out std_logic;                                        -- of_wr
			of_wrfull          : in  std_logic                     := 'X';             -- of_wrfull
			if_d               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- if_d
			if_rd              : out std_logic;                                        -- if_rd
			if_rdempty         : in  std_logic                     := 'X';             -- if_rdempty
			fifo_rst           : out std_logic                                         -- fifo_rst
		);
	end component avs_fifo_int;

	component factory_bridge_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			avalon_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avalon_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			avalon_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			avalon_read        : out std_logic;                                        -- read
			avalon_write       : out std_logic;                                        -- write
			avalon_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			avalon_address     : out std_logic_vector(20 downto 0);                    -- address
			address            : in  std_logic_vector(20 downto 0) := (others => 'X'); -- export
			byte_enable        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			read               : in  std_logic                     := 'X';             -- export
			write              : in  std_logic                     := 'X';             -- export
			write_data         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			acknowledge        : out std_logic;                                        -- export
			read_data          : out std_logic_vector(31 downto 0)                     -- export
		);
	end component factory_bridge_0;

	component altera_dual_boot is
		generic (
			INTENDED_DEVICE_FAMILY : string  := "";
			CONFIG_CYCLE           : integer := 28;
			RESET_TIMER_CYCLE      : integer := 40
		);
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			nreset             : in  std_logic                     := 'X';             -- reset_n
			avmm_rcv_address   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avmm_rcv_read      : in  std_logic                     := 'X';             -- read
			avmm_rcv_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_rcv_write     : in  std_logic                     := 'X';             -- write
			avmm_rcv_readdata  : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component altera_dual_boot;

	component i2c_opencores is
		port (
			wb_clk_i   : in    std_logic                    := 'X';             -- clk
			wb_rst_i   : in    std_logic                    := 'X';             -- reset
			scl_pad_io : inout std_logic                    := 'X';             -- export
			sda_pad_io : inout std_logic                    := 'X';             -- export
			wb_adr_i   : in    std_logic_vector(2 downto 0) := (others => 'X'); -- address
			wb_dat_i   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			wb_dat_o   : out   std_logic_vector(7 downto 0);                    -- readdata
			wb_we_i    : in    std_logic                    := 'X';             -- write
			wb_stb_i   : in    std_logic                    := 'X';             -- chipselect
			wb_ack_o   : out   std_logic;                                       -- waitrequest_n
			wb_inta_o  : out   std_logic                                        -- irq
		);
	end component i2c_opencores;

	component altera_onchip_flash is
		generic (
			INIT_FILENAME                       : string  := "";
			INIT_FILENAME_SIM                   : string  := "";
			DEVICE_FAMILY                       : string  := "Unknown";
			PART_NAME                           : string  := "Unknown";
			DEVICE_ID                           : string  := "Unknown";
			SECTOR1_START_ADDR                  : integer := 0;
			SECTOR1_END_ADDR                    : integer := 0;
			SECTOR2_START_ADDR                  : integer := 0;
			SECTOR2_END_ADDR                    : integer := 0;
			SECTOR3_START_ADDR                  : integer := 0;
			SECTOR3_END_ADDR                    : integer := 0;
			SECTOR4_START_ADDR                  : integer := 0;
			SECTOR4_END_ADDR                    : integer := 0;
			SECTOR5_START_ADDR                  : integer := 0;
			SECTOR5_END_ADDR                    : integer := 0;
			MIN_VALID_ADDR                      : integer := 0;
			MAX_VALID_ADDR                      : integer := 0;
			MIN_UFM_VALID_ADDR                  : integer := 0;
			MAX_UFM_VALID_ADDR                  : integer := 0;
			SECTOR1_MAP                         : integer := 0;
			SECTOR2_MAP                         : integer := 0;
			SECTOR3_MAP                         : integer := 0;
			SECTOR4_MAP                         : integer := 0;
			SECTOR5_MAP                         : integer := 0;
			ADDR_RANGE1_END_ADDR                : integer := 0;
			ADDR_RANGE2_END_ADDR                : integer := 0;
			ADDR_RANGE1_OFFSET                  : integer := 0;
			ADDR_RANGE2_OFFSET                  : integer := 0;
			ADDR_RANGE3_OFFSET                  : integer := 0;
			AVMM_DATA_ADDR_WIDTH                : integer := 19;
			AVMM_DATA_DATA_WIDTH                : integer := 32;
			AVMM_DATA_BURSTCOUNT_WIDTH          : integer := 4;
			SECTOR_READ_PROTECTION_MODE         : integer := 31;
			FLASH_SEQ_READ_DATA_COUNT           : integer := 2;
			FLASH_ADDR_ALIGNMENT_BITS           : integer := 1;
			FLASH_READ_CYCLE_MAX_INDEX          : integer := 4;
			FLASH_RESET_CYCLE_MAX_INDEX         : integer := 29;
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  : integer := 112;
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX : integer := 40603248;
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX : integer := 35382;
			PARALLEL_MODE                       : boolean := true;
			READ_AND_WRITE_MODE                 : boolean := true;
			WRAPPING_BURST_MODE                 : boolean := false;
			IS_DUAL_BOOT                        : string  := "False";
			IS_ERAM_SKIP                        : string  := "False";
			IS_COMPRESSED_IMAGE                 : string  := "False"
		);
		port (
			clock                   : in  std_logic                     := 'X';             -- clk
			reset_n                 : in  std_logic                     := 'X';             -- reset_n
			avmm_data_addr          : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			avmm_data_read          : in  std_logic                     := 'X';             -- read
			avmm_data_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_data_write         : in  std_logic                     := 'X';             -- write
			avmm_data_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avmm_data_waitrequest   : out std_logic;                                        -- waitrequest
			avmm_data_readdatavalid : out std_logic;                                        -- readdatavalid
			avmm_data_burstcount    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			avmm_csr_addr           : in  std_logic                     := 'X';             -- address
			avmm_csr_read           : in  std_logic                     := 'X';             -- read
			avmm_csr_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_csr_write          : in  std_logic                     := 'X';             -- write
			avmm_csr_readdata       : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component altera_onchip_flash;

	component factory_pio_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component factory_pio_0;

	component factory_mm_interconnect_0 is
		port (
			clk_0_clk_clk                              : in  std_logic                     := 'X';             -- clk
			bridge_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			bridge_0_avalon_master_address             : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			bridge_0_avalon_master_waitrequest         : out std_logic;                                        -- waitrequest
			bridge_0_avalon_master_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			bridge_0_avalon_master_read                : in  std_logic                     := 'X';             -- read
			bridge_0_avalon_master_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			bridge_0_avalon_master_write               : in  std_logic                     := 'X';             -- write
			bridge_0_avalon_master_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_fifo_int_0_avs_s0_address              : out std_logic_vector(7 downto 0);                     -- address
			avs_fifo_int_0_avs_s0_write                : out std_logic;                                        -- write
			avs_fifo_int_0_avs_s0_read                 : out std_logic;                                        -- read
			avs_fifo_int_0_avs_s0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avs_fifo_int_0_avs_s0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			avs_fifo_int_0_avs_s0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			dual_boot_0_avalon_address                 : out std_logic_vector(2 downto 0);                     -- address
			dual_boot_0_avalon_write                   : out std_logic;                                        -- write
			dual_boot_0_avalon_read                    : out std_logic;                                        -- read
			dual_boot_0_avalon_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dual_boot_0_avalon_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			i2c_opencores_0_avalon_slave_0_address     : out std_logic_vector(2 downto 0);                     -- address
			i2c_opencores_0_avalon_slave_0_write       : out std_logic;                                        -- write
			i2c_opencores_0_avalon_slave_0_readdata    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_opencores_0_avalon_slave_0_writedata   : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_opencores_0_avalon_slave_0_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			i2c_opencores_0_avalon_slave_0_chipselect  : out std_logic;                                        -- chipselect
			onchip_flash_0_csr_address                 : out std_logic_vector(0 downto 0);                     -- address
			onchip_flash_0_csr_write                   : out std_logic;                                        -- write
			onchip_flash_0_csr_read                    : out std_logic;                                        -- read
			onchip_flash_0_csr_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_flash_0_csr_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_flash_0_data_address                : out std_logic_vector(17 downto 0);                    -- address
			onchip_flash_0_data_write                  : out std_logic;                                        -- write
			onchip_flash_0_data_read                   : out std_logic;                                        -- read
			onchip_flash_0_data_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_flash_0_data_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_flash_0_data_burstcount             : out std_logic_vector(3 downto 0);                     -- burstcount
			onchip_flash_0_data_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			onchip_flash_0_data_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			pio_0_s1_address                           : out std_logic_vector(2 downto 0);                     -- address
			pio_0_s1_write                             : out std_logic;                                        -- write
			pio_0_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_0_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			pio_0_s1_chipselect                        : out std_logic                                         -- chipselect
		);
	end component factory_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal bridge_0_avalon_master_readdata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:bridge_0_avalon_master_readdata -> bridge_0:avalon_readdata
	signal bridge_0_avalon_master_waitrequest                          : std_logic;                     -- mm_interconnect_0:bridge_0_avalon_master_waitrequest -> bridge_0:avalon_waitrequest
	signal bridge_0_avalon_master_byteenable                           : std_logic_vector(3 downto 0);  -- bridge_0:avalon_byteenable -> mm_interconnect_0:bridge_0_avalon_master_byteenable
	signal bridge_0_avalon_master_read                                 : std_logic;                     -- bridge_0:avalon_read -> mm_interconnect_0:bridge_0_avalon_master_read
	signal bridge_0_avalon_master_address                              : std_logic_vector(20 downto 0); -- bridge_0:avalon_address -> mm_interconnect_0:bridge_0_avalon_master_address
	signal bridge_0_avalon_master_write                                : std_logic;                     -- bridge_0:avalon_write -> mm_interconnect_0:bridge_0_avalon_master_write
	signal bridge_0_avalon_master_writedata                            : std_logic_vector(31 downto 0); -- bridge_0:avalon_writedata -> mm_interconnect_0:bridge_0_avalon_master_writedata
	signal mm_interconnect_0_dual_boot_0_avalon_readdata               : std_logic_vector(31 downto 0); -- dual_boot_0:avmm_rcv_readdata -> mm_interconnect_0:dual_boot_0_avalon_readdata
	signal mm_interconnect_0_dual_boot_0_avalon_address                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:dual_boot_0_avalon_address -> dual_boot_0:avmm_rcv_address
	signal mm_interconnect_0_dual_boot_0_avalon_read                   : std_logic;                     -- mm_interconnect_0:dual_boot_0_avalon_read -> dual_boot_0:avmm_rcv_read
	signal mm_interconnect_0_dual_boot_0_avalon_write                  : std_logic;                     -- mm_interconnect_0:dual_boot_0_avalon_write -> dual_boot_0:avmm_rcv_write
	signal mm_interconnect_0_dual_boot_0_avalon_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:dual_boot_0_avalon_writedata -> dual_boot_0:avmm_rcv_writedata
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect : std_logic;                     -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_chipselect -> i2c_opencores_0:wb_stb_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata   : std_logic_vector(7 downto 0);  -- i2c_opencores_0:wb_dat_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_readdata
	signal i2c_opencores_0_avalon_slave_0_waitrequest                  : std_logic;                     -- i2c_opencores_0:wb_ack_o -> i2c_opencores_0_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_address -> i2c_opencores_0:wb_adr_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write      : std_logic;                     -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_write -> i2c_opencores_0:wb_we_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_writedata -> i2c_opencores_0:wb_dat_i
	signal mm_interconnect_0_avs_fifo_int_0_avs_s0_readdata            : std_logic_vector(31 downto 0); -- avs_fifo_int_0:avs_s0_readdata -> mm_interconnect_0:avs_fifo_int_0_avs_s0_readdata
	signal mm_interconnect_0_avs_fifo_int_0_avs_s0_waitrequest         : std_logic;                     -- avs_fifo_int_0:avs_s0_waitrequest -> mm_interconnect_0:avs_fifo_int_0_avs_s0_waitrequest
	signal mm_interconnect_0_avs_fifo_int_0_avs_s0_address             : std_logic_vector(7 downto 0);  -- mm_interconnect_0:avs_fifo_int_0_avs_s0_address -> avs_fifo_int_0:avs_s0_address
	signal mm_interconnect_0_avs_fifo_int_0_avs_s0_read                : std_logic;                     -- mm_interconnect_0:avs_fifo_int_0_avs_s0_read -> avs_fifo_int_0:avs_s0_read
	signal mm_interconnect_0_avs_fifo_int_0_avs_s0_write               : std_logic;                     -- mm_interconnect_0:avs_fifo_int_0_avs_s0_write -> avs_fifo_int_0:avs_s0_write
	signal mm_interconnect_0_avs_fifo_int_0_avs_s0_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:avs_fifo_int_0_avs_s0_writedata -> avs_fifo_int_0:avs_s0_writedata
	signal mm_interconnect_0_onchip_flash_0_csr_readdata               : std_logic_vector(31 downto 0); -- onchip_flash_0:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_0_csr_readdata
	signal mm_interconnect_0_onchip_flash_0_csr_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	signal mm_interconnect_0_onchip_flash_0_csr_read                   : std_logic;                     -- mm_interconnect_0:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	signal mm_interconnect_0_onchip_flash_0_csr_write                  : std_logic;                     -- mm_interconnect_0:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	signal mm_interconnect_0_onchip_flash_0_csr_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	signal mm_interconnect_0_onchip_flash_0_data_readdata              : std_logic_vector(31 downto 0); -- onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	signal mm_interconnect_0_onchip_flash_0_data_waitrequest           : std_logic;                     -- onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	signal mm_interconnect_0_onchip_flash_0_data_address               : std_logic_vector(17 downto 0); -- mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	signal mm_interconnect_0_onchip_flash_0_data_read                  : std_logic;                     -- mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	signal mm_interconnect_0_onchip_flash_0_data_readdatavalid         : std_logic;                     -- onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	signal mm_interconnect_0_onchip_flash_0_data_write                 : std_logic;                     -- mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	signal mm_interconnect_0_onchip_flash_0_data_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	signal mm_interconnect_0_onchip_flash_0_data_burstcount            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	signal mm_interconnect_0_pio_0_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	signal mm_interconnect_0_pio_0_s1_readdata                         : std_logic_vector(31 downto 0); -- pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	signal mm_interconnect_0_pio_0_s1_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:pio_0_s1_address -> pio_0:address
	signal mm_interconnect_0_pio_0_s1_write                            : std_logic;                     -- mm_interconnect_0:pio_0_s1_write -> mm_interconnect_0_pio_0_s1_write:in
	signal mm_interconnect_0_pio_0_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	signal rst_controller_reset_out_reset                              : std_logic;                     -- rst_controller:reset_out -> [avs_fifo_int_0:reset_reset, bridge_0:reset, i2c_opencores_0:wb_rst_i, mm_interconnect_0:bridge_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                     : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv        : std_logic;                     -- i2c_opencores_0_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_pio_0_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_pio_0_s1_write:inv -> pio_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_reset_out_reset:inv -> [dual_boot_0:nreset, onchip_flash_0:reset_n, pio_0:reset_n]

begin

	avs_fifo_int_0 : component avs_fifo_int
		port map (
			avs_s0_address     => mm_interconnect_0_avs_fifo_int_0_avs_s0_address,     -- avs_s0.address
			avs_s0_read        => mm_interconnect_0_avs_fifo_int_0_avs_s0_read,        --       .read
			avs_s0_readdata    => mm_interconnect_0_avs_fifo_int_0_avs_s0_readdata,    --       .readdata
			avs_s0_write       => mm_interconnect_0_avs_fifo_int_0_avs_s0_write,       --       .write
			avs_s0_writedata   => mm_interconnect_0_avs_fifo_int_0_avs_s0_writedata,   --       .writedata
			avs_s0_waitrequest => mm_interconnect_0_avs_fifo_int_0_avs_s0_waitrequest, --       .waitrequest
			clock_clk          => clk_clk,                                             --  clock.clk
			reset_reset        => rst_controller_reset_out_reset,                      --  reset.reset
			of_d               => extfifo_of_d,                                        --    coe.of_d
			of_wr              => extfifo_of_wr,                                       --       .of_wr
			of_wrfull          => extfifo_of_wrfull,                                   --       .of_wrfull
			if_d               => extfifo_if_d,                                        --       .if_d
			if_rd              => extfifo_if_rd,                                       --       .if_rd
			if_rdempty         => extfifo_if_rdempty,                                  --       .if_rdempty
			fifo_rst           => extfifo_fifo_rst                                     --       .fifo_rst
		);

	bridge_0 : component factory_bridge_0
		port map (
			clk                => clk_clk,                            --                clk.clk
			reset              => rst_controller_reset_out_reset,     --              reset.reset
			avalon_readdata    => bridge_0_avalon_master_readdata,    --      avalon_master.readdata
			avalon_waitrequest => bridge_0_avalon_master_waitrequest, --                   .waitrequest
			avalon_byteenable  => bridge_0_avalon_master_byteenable,  --                   .byteenable
			avalon_read        => bridge_0_avalon_master_read,        --                   .read
			avalon_write       => bridge_0_avalon_master_write,       --                   .write
			avalon_writedata   => bridge_0_avalon_master_writedata,   --                   .writedata
			avalon_address     => bridge_0_avalon_master_address,     --                   .address
			address            => bridge_0_address,                   -- external_interface.export
			byte_enable        => bridge_0_byte_enable,               --                   .export
			read               => bridge_0_read,                      --                   .export
			write              => bridge_0_write,                     --                   .export
			write_data         => bridge_0_write_data,                --                   .export
			acknowledge        => bridge_0_acknowledge,               --                   .export
			read_data          => bridge_0_read_data                  --                   .export
		);

	dual_boot_0 : component altera_dual_boot
		generic map (
			INTENDED_DEVICE_FAMILY => "MAX 10",
			CONFIG_CYCLE           => 15,
			RESET_TIMER_CYCLE      => 21
		)
		port map (
			clk                => clk_clk,                                        --    clk.clk
			nreset             => rst_controller_reset_out_reset_ports_inv,       -- nreset.reset_n
			avmm_rcv_address   => mm_interconnect_0_dual_boot_0_avalon_address,   -- avalon.address
			avmm_rcv_read      => mm_interconnect_0_dual_boot_0_avalon_read,      --       .read
			avmm_rcv_writedata => mm_interconnect_0_dual_boot_0_avalon_writedata, --       .writedata
			avmm_rcv_write     => mm_interconnect_0_dual_boot_0_avalon_write,     --       .write
			avmm_rcv_readdata  => mm_interconnect_0_dual_boot_0_avalon_readdata   --       .readdata
		);

	i2c_opencores_0 : component i2c_opencores
		port map (
			wb_clk_i   => clk_clk,                                                     --            clock.clk
			wb_rst_i   => rst_controller_reset_out_reset,                              --      clock_reset.reset
			scl_pad_io => scl_export,                                                  --       export_scl.export
			sda_pad_io => sda_export,                                                  --       export_sda.export
			wb_adr_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_opencores_0_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			wb_inta_o  => open                                                         -- interrupt_sender.irq
		);

	onchip_flash_0 : component altera_onchip_flash
		generic map (
			INIT_FILENAME                       => "",
			INIT_FILENAME_SIM                   => "",
			DEVICE_FAMILY                       => "MAX 10",
			PART_NAME                           => "10M16SAU169I7G",
			DEVICE_ID                           => "16",
			SECTOR1_START_ADDR                  => 0,
			SECTOR1_END_ADDR                    => 4095,
			SECTOR2_START_ADDR                  => 4096,
			SECTOR2_END_ADDR                    => 8191,
			SECTOR3_START_ADDR                  => 8192,
			SECTOR3_END_ADDR                    => 47103,
			SECTOR4_START_ADDR                  => 47104,
			SECTOR4_END_ADDR                    => 75775,
			SECTOR5_START_ADDR                  => 75776,
			SECTOR5_END_ADDR                    => 143359,
			MIN_VALID_ADDR                      => 0,
			MAX_VALID_ADDR                      => 143359,
			MIN_UFM_VALID_ADDR                  => 0,
			MAX_UFM_VALID_ADDR                  => 8191,
			SECTOR1_MAP                         => 1,
			SECTOR2_MAP                         => 2,
			SECTOR3_MAP                         => 3,
			SECTOR4_MAP                         => 4,
			SECTOR5_MAP                         => 5,
			ADDR_RANGE1_END_ADDR                => 143359,
			ADDR_RANGE2_END_ADDR                => 143359,
			ADDR_RANGE1_OFFSET                  => 1024,
			ADDR_RANGE2_OFFSET                  => 0,
			ADDR_RANGE3_OFFSET                  => 0,
			AVMM_DATA_ADDR_WIDTH                => 18,
			AVMM_DATA_DATA_WIDTH                => 32,
			AVMM_DATA_BURSTCOUNT_WIDTH          => 4,
			SECTOR_READ_PROTECTION_MODE         => 0,
			FLASH_SEQ_READ_DATA_COUNT           => 4,
			FLASH_ADDR_ALIGNMENT_BITS           => 2,
			FLASH_READ_CYCLE_MAX_INDEX          => 4,
			FLASH_RESET_CYCLE_MAX_INDEX         => 7,
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  => 36,
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX => 10752027,
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX => 9369,
			PARALLEL_MODE                       => true,
			READ_AND_WRITE_MODE                 => true,
			WRAPPING_BURST_MODE                 => false,
			IS_DUAL_BOOT                        => "True",
			IS_ERAM_SKIP                        => "True",
			IS_COMPRESSED_IMAGE                 => "True"
		)
		port map (
			clock                   => clk_clk,                                             --    clk.clk
			reset_n                 => rst_controller_reset_out_reset_ports_inv,            -- nreset.reset_n
			avmm_data_addr          => mm_interconnect_0_onchip_flash_0_data_address,       --   data.address
			avmm_data_read          => mm_interconnect_0_onchip_flash_0_data_read,          --       .read
			avmm_data_writedata     => mm_interconnect_0_onchip_flash_0_data_writedata,     --       .writedata
			avmm_data_write         => mm_interconnect_0_onchip_flash_0_data_write,         --       .write
			avmm_data_readdata      => mm_interconnect_0_onchip_flash_0_data_readdata,      --       .readdata
			avmm_data_waitrequest   => mm_interconnect_0_onchip_flash_0_data_waitrequest,   --       .waitrequest
			avmm_data_readdatavalid => mm_interconnect_0_onchip_flash_0_data_readdatavalid, --       .readdatavalid
			avmm_data_burstcount    => mm_interconnect_0_onchip_flash_0_data_burstcount,    --       .burstcount
			avmm_csr_addr           => mm_interconnect_0_onchip_flash_0_csr_address(0),     --    csr.address
			avmm_csr_read           => mm_interconnect_0_onchip_flash_0_csr_read,           --       .read
			avmm_csr_writedata      => mm_interconnect_0_onchip_flash_0_csr_writedata,      --       .writedata
			avmm_csr_write          => mm_interconnect_0_onchip_flash_0_csr_write,          --       .write
			avmm_csr_readdata       => mm_interconnect_0_onchip_flash_0_csr_readdata        --       .readdata
		);

	pio_0 : component factory_pio_0
		port map (
			clk        => clk_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pio_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_0_s1_readdata,        --                    .readdata
			out_port   => pio_0_export                                -- external_connection.export
		);

	mm_interconnect_0 : component factory_mm_interconnect_0
		port map (
			clk_0_clk_clk                              => clk_clk,                                                     --                            clk_0_clk.clk
			bridge_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- bridge_0_reset_reset_bridge_in_reset.reset
			bridge_0_avalon_master_address             => bridge_0_avalon_master_address,                              --               bridge_0_avalon_master.address
			bridge_0_avalon_master_waitrequest         => bridge_0_avalon_master_waitrequest,                          --                                     .waitrequest
			bridge_0_avalon_master_byteenable          => bridge_0_avalon_master_byteenable,                           --                                     .byteenable
			bridge_0_avalon_master_read                => bridge_0_avalon_master_read,                                 --                                     .read
			bridge_0_avalon_master_readdata            => bridge_0_avalon_master_readdata,                             --                                     .readdata
			bridge_0_avalon_master_write               => bridge_0_avalon_master_write,                                --                                     .write
			bridge_0_avalon_master_writedata           => bridge_0_avalon_master_writedata,                            --                                     .writedata
			avs_fifo_int_0_avs_s0_address              => mm_interconnect_0_avs_fifo_int_0_avs_s0_address,             --                avs_fifo_int_0_avs_s0.address
			avs_fifo_int_0_avs_s0_write                => mm_interconnect_0_avs_fifo_int_0_avs_s0_write,               --                                     .write
			avs_fifo_int_0_avs_s0_read                 => mm_interconnect_0_avs_fifo_int_0_avs_s0_read,                --                                     .read
			avs_fifo_int_0_avs_s0_readdata             => mm_interconnect_0_avs_fifo_int_0_avs_s0_readdata,            --                                     .readdata
			avs_fifo_int_0_avs_s0_writedata            => mm_interconnect_0_avs_fifo_int_0_avs_s0_writedata,           --                                     .writedata
			avs_fifo_int_0_avs_s0_waitrequest          => mm_interconnect_0_avs_fifo_int_0_avs_s0_waitrequest,         --                                     .waitrequest
			dual_boot_0_avalon_address                 => mm_interconnect_0_dual_boot_0_avalon_address,                --                   dual_boot_0_avalon.address
			dual_boot_0_avalon_write                   => mm_interconnect_0_dual_boot_0_avalon_write,                  --                                     .write
			dual_boot_0_avalon_read                    => mm_interconnect_0_dual_boot_0_avalon_read,                   --                                     .read
			dual_boot_0_avalon_readdata                => mm_interconnect_0_dual_boot_0_avalon_readdata,               --                                     .readdata
			dual_boot_0_avalon_writedata               => mm_interconnect_0_dual_boot_0_avalon_writedata,              --                                     .writedata
			i2c_opencores_0_avalon_slave_0_address     => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address,    --       i2c_opencores_0_avalon_slave_0.address
			i2c_opencores_0_avalon_slave_0_write       => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write,      --                                     .write
			i2c_opencores_0_avalon_slave_0_readdata    => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata,   --                                     .readdata
			i2c_opencores_0_avalon_slave_0_writedata   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata,  --                                     .writedata
			i2c_opencores_0_avalon_slave_0_waitrequest => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv,        --                                     .waitrequest
			i2c_opencores_0_avalon_slave_0_chipselect  => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect, --                                     .chipselect
			onchip_flash_0_csr_address                 => mm_interconnect_0_onchip_flash_0_csr_address,                --                   onchip_flash_0_csr.address
			onchip_flash_0_csr_write                   => mm_interconnect_0_onchip_flash_0_csr_write,                  --                                     .write
			onchip_flash_0_csr_read                    => mm_interconnect_0_onchip_flash_0_csr_read,                   --                                     .read
			onchip_flash_0_csr_readdata                => mm_interconnect_0_onchip_flash_0_csr_readdata,               --                                     .readdata
			onchip_flash_0_csr_writedata               => mm_interconnect_0_onchip_flash_0_csr_writedata,              --                                     .writedata
			onchip_flash_0_data_address                => mm_interconnect_0_onchip_flash_0_data_address,               --                  onchip_flash_0_data.address
			onchip_flash_0_data_write                  => mm_interconnect_0_onchip_flash_0_data_write,                 --                                     .write
			onchip_flash_0_data_read                   => mm_interconnect_0_onchip_flash_0_data_read,                  --                                     .read
			onchip_flash_0_data_readdata               => mm_interconnect_0_onchip_flash_0_data_readdata,              --                                     .readdata
			onchip_flash_0_data_writedata              => mm_interconnect_0_onchip_flash_0_data_writedata,             --                                     .writedata
			onchip_flash_0_data_burstcount             => mm_interconnect_0_onchip_flash_0_data_burstcount,            --                                     .burstcount
			onchip_flash_0_data_readdatavalid          => mm_interconnect_0_onchip_flash_0_data_readdatavalid,         --                                     .readdatavalid
			onchip_flash_0_data_waitrequest            => mm_interconnect_0_onchip_flash_0_data_waitrequest,           --                                     .waitrequest
			pio_0_s1_address                           => mm_interconnect_0_pio_0_s1_address,                          --                             pio_0_s1.address
			pio_0_s1_write                             => mm_interconnect_0_pio_0_s1_write,                            --                                     .write
			pio_0_s1_readdata                          => mm_interconnect_0_pio_0_s1_readdata,                         --                                     .readdata
			pio_0_s1_writedata                         => mm_interconnect_0_pio_0_s1_writedata,                        --                                     .writedata
			pio_0_s1_chipselect                        => mm_interconnect_0_pio_0_s1_chipselect                        --                                     .chipselect
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv <= not i2c_opencores_0_avalon_slave_0_waitrequest;

	mm_interconnect_0_pio_0_s1_write_ports_inv <= not mm_interconnect_0_pio_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of factory
