-- lms_ctr.vhd

-- Generated using ACDS version 18.0 614

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity lms_ctr is
	port (
		avm_m0_address                          : out   std_logic_vector(7 downto 0);                     --                           avm_m0.address
		avm_m0_read                             : out   std_logic;                                        --                                 .read
		avm_m0_waitrequest                      : in    std_logic                     := '0';             --                                 .waitrequest
		avm_m0_readdata                         : in    std_logic_vector(7 downto 0)  := (others => '0'); --                                 .readdata
		avm_m0_write                            : out   std_logic;                                        --                                 .write
		avm_m0_writedata                        : out   std_logic_vector(7 downto 0);                     --                                 .writedata
		avm_m0_readdatavalid                    : in    std_logic                     := '0';             --                                 .readdatavalid
		avm_m0_clk_clk                          : out   std_logic;                                        --                       avm_m0_clk.clk
		avm_m0_reset_reset                      : out   std_logic;                                        --                     avm_m0_reset.reset
		clk_clk                                 : in    std_logic                     := '0';             --                              clk.clk
		dac_spi_ext_MISO                        : in    std_logic                     := '0';             --                      dac_spi_ext.MISO
		dac_spi_ext_MOSI                        : out   std_logic;                                        --                                 .MOSI
		dac_spi_ext_SCLK                        : out   std_logic;                                        --                                 .SCLK
		dac_spi_ext_SS_n                        : out   std_logic;                                        --                                 .SS_n
		exfifo_if_d_export                      : in    std_logic_vector(31 downto 0) := (others => '0'); --                      exfifo_if_d.export
		exfifo_if_rd_export                     : out   std_logic;                                        --                     exfifo_if_rd.export
		exfifo_if_rdempty_export                : in    std_logic                     := '0';             --                exfifo_if_rdempty.export
		exfifo_of_d_export                      : out   std_logic_vector(31 downto 0);                    --                      exfifo_of_d.export
		exfifo_of_wr_export                     : out   std_logic;                                        --                     exfifo_of_wr.export
		exfifo_of_wrfull_export                 : in    std_logic                     := '0';             --                 exfifo_of_wrfull.export
		exfifo_rst_export                       : out   std_logic;                                        --                       exfifo_rst.export
		flash_spi_MISO                          : in    std_logic                     := '0';             --                        flash_spi.MISO
		flash_spi_MOSI                          : out   std_logic;                                        --                                 .MOSI
		flash_spi_SCLK                          : out   std_logic;                                        --                                 .SCLK
		flash_spi_SS_n                          : out   std_logic;                                        --                                 .SS_n
		fpga_spi_ext_MISO                       : in    std_logic                     := '0';             --                     fpga_spi_ext.MISO
		fpga_spi_ext_MOSI                       : out   std_logic;                                        --                                 .MOSI
		fpga_spi_ext_SCLK                       : out   std_logic;                                        --                                 .SCLK
		fpga_spi_ext_SS_n                       : out   std_logic_vector(2 downto 0);                     --                                 .SS_n
		i2c_scl_export                          : inout std_logic                     := '0';             --                          i2c_scl.export
		i2c_sda_export                          : inout std_logic                     := '0';             --                          i2c_sda.export
		leds_external_connection_export         : out   std_logic_vector(7 downto 0);                     --         leds_external_connection.export
		lms_ctr_gpio_external_connection_export : out   std_logic_vector(3 downto 0);                     -- lms_ctr_gpio_external_connection.export
		reset_reset_n                           : in    std_logic                     := '0';             --                            reset.reset_n
		switch_external_connection_export       : in    std_logic_vector(7 downto 0)  := (others => '0'); --       switch_external_connection.export
		vctcxo_tamer_0_ctrl_export              : in    std_logic_vector(3 downto 0)  := (others => '0')  --              vctcxo_tamer_0_ctrl.export
	);
end entity lms_ctr;

architecture rtl of lms_ctr is
	component avfifo is
		generic (
			width : integer := 32
		);
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			chipselect     : in  std_logic                     := 'X';             -- chipselect
			write          : in  std_logic                     := 'X';             -- write
			writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			read           : in  std_logic                     := 'X';             -- read
			readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			rsi_nrst       : in  std_logic                     := 'X';             -- reset_n
			coe_if_d       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			coe_if_rd      : out std_logic;                                        -- export
			coe_of_wrfull  : in  std_logic                     := 'X';             -- export
			coe_of_wr      : out std_logic;                                        -- export
			coe_of_d       : out std_logic_vector(31 downto 0);                    -- export
			coe_if_rdempty : in  std_logic                     := 'X';             -- export
			coe_fifo_rst   : out std_logic                                         -- export
		);
	end component avfifo;

	component Avalon_MM_external is
		port (
			avs_s0_address       : in  std_logic_vector(7 downto 0) := (others => 'X'); -- address
			avs_s0_read          : in  std_logic                    := 'X';             -- read
			avs_s0_readdata      : out std_logic_vector(7 downto 0);                    -- readdata
			avs_s0_write         : in  std_logic                    := 'X';             -- write
			avs_s0_writedata     : in  std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			avs_s0_waitrequest   : out std_logic;                                       -- waitrequest
			avs_s0_readdatavalid : out std_logic;                                       -- readdatavalid
			clock_clk            : in  std_logic                    := 'X';             -- clk
			reset_reset          : in  std_logic                    := 'X';             -- reset
			avm_m0_address       : out std_logic_vector(7 downto 0);                    -- address
			avm_m0_read          : out std_logic;                                       -- read
			avm_m0_waitrequest   : in  std_logic                    := 'X';             -- waitrequest
			avm_m0_readdata      : in  std_logic_vector(7 downto 0) := (others => 'X'); -- readdata
			avm_m0_write         : out std_logic;                                       -- write
			avm_m0_writedata     : out std_logic_vector(7 downto 0);                    -- writedata
			avm_m0_readdatavalid : in  std_logic                    := 'X';             -- readdatavalid
			clock_source_clk     : out std_logic;                                       -- clk
			reset_source_reset   : out std_logic                                        -- reset
		);
	end component Avalon_MM_external;

	component lms_ctr_dac_spi is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component lms_ctr_dac_spi;

	component altera_dual_boot is
		generic (
			INTENDED_DEVICE_FAMILY : string  := "";
			CONFIG_CYCLE           : integer := 28;
			RESET_TIMER_CYCLE      : integer := 40
		);
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			nreset             : in  std_logic                     := 'X';             -- reset_n
			avmm_rcv_address   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avmm_rcv_read      : in  std_logic                     := 'X';             -- read
			avmm_rcv_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_rcv_write     : in  std_logic                     := 'X';             -- write
			avmm_rcv_readdata  : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component altera_dual_boot;

	component lms_ctr_flash_spi is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component lms_ctr_flash_spi;

	component lms_ctr_fpga_spi is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic_vector(2 downto 0)                      -- export
		);
	end component lms_ctr_fpga_spi;

	component i2c_opencores is
		port (
			wb_clk_i   : in    std_logic                    := 'X';             -- clk
			wb_rst_i   : in    std_logic                    := 'X';             -- reset
			scl_pad_io : inout std_logic                    := 'X';             -- export
			sda_pad_io : inout std_logic                    := 'X';             -- export
			wb_adr_i   : in    std_logic_vector(2 downto 0) := (others => 'X'); -- address
			wb_dat_i   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			wb_dat_o   : out   std_logic_vector(7 downto 0);                    -- readdata
			wb_we_i    : in    std_logic                    := 'X';             -- write
			wb_stb_i   : in    std_logic                    := 'X';             -- chipselect
			wb_ack_o   : out   std_logic;                                       -- waitrequest_n
			wb_inta_o  : out   std_logic                                        -- irq
		);
	end component i2c_opencores;

	component lms_ctr_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component lms_ctr_leds;

	component lms_ctr_lms_ctr_gpio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component lms_ctr_lms_ctr_gpio;

	component lms_ctr_nios2_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(21 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(21 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			E_ci_result                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			D_ci_a                              : out std_logic_vector(4 downto 0);                     -- a
			D_ci_b                              : out std_logic_vector(4 downto 0);                     -- b
			D_ci_c                              : out std_logic_vector(4 downto 0);                     -- c
			D_ci_n                              : out std_logic_vector(7 downto 0);                     -- n
			D_ci_readra                         : out std_logic;                                        -- readra
			D_ci_readrb                         : out std_logic;                                        -- readrb
			D_ci_writerc                        : out std_logic;                                        -- writerc
			E_ci_dataa                          : out std_logic_vector(31 downto 0);                    -- dataa
			E_ci_datab                          : out std_logic_vector(31 downto 0);                    -- datab
			E_ci_multi_clock                    : out std_logic;                                        -- clk
			E_ci_multi_reset                    : out std_logic;                                        -- reset
			E_ci_multi_reset_req                : out std_logic;                                        -- reset_req
			W_ci_estatus                        : out std_logic;                                        -- estatus
			W_ci_ipending                       : out std_logic_vector(31 downto 0)                     -- ipending
		);
	end component lms_ctr_nios2_cpu;

	component bitswap_qsys is
		port (
			dataa  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			datab  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			result : out std_logic_vector(31 downto 0)                     -- result
		);
	end component bitswap_qsys;

	component altera_onchip_flash is
		generic (
			INIT_FILENAME                       : string  := "";
			INIT_FILENAME_SIM                   : string  := "";
			DEVICE_FAMILY                       : string  := "Unknown";
			PART_NAME                           : string  := "Unknown";
			DEVICE_ID                           : string  := "Unknown";
			SECTOR1_START_ADDR                  : integer := 0;
			SECTOR1_END_ADDR                    : integer := 0;
			SECTOR2_START_ADDR                  : integer := 0;
			SECTOR2_END_ADDR                    : integer := 0;
			SECTOR3_START_ADDR                  : integer := 0;
			SECTOR3_END_ADDR                    : integer := 0;
			SECTOR4_START_ADDR                  : integer := 0;
			SECTOR4_END_ADDR                    : integer := 0;
			SECTOR5_START_ADDR                  : integer := 0;
			SECTOR5_END_ADDR                    : integer := 0;
			MIN_VALID_ADDR                      : integer := 0;
			MAX_VALID_ADDR                      : integer := 0;
			MIN_UFM_VALID_ADDR                  : integer := 0;
			MAX_UFM_VALID_ADDR                  : integer := 0;
			SECTOR1_MAP                         : integer := 0;
			SECTOR2_MAP                         : integer := 0;
			SECTOR3_MAP                         : integer := 0;
			SECTOR4_MAP                         : integer := 0;
			SECTOR5_MAP                         : integer := 0;
			ADDR_RANGE1_END_ADDR                : integer := 0;
			ADDR_RANGE2_END_ADDR                : integer := 0;
			ADDR_RANGE1_OFFSET                  : integer := 0;
			ADDR_RANGE2_OFFSET                  : integer := 0;
			ADDR_RANGE3_OFFSET                  : integer := 0;
			AVMM_DATA_ADDR_WIDTH                : integer := 19;
			AVMM_DATA_DATA_WIDTH                : integer := 32;
			AVMM_DATA_BURSTCOUNT_WIDTH          : integer := 4;
			SECTOR_READ_PROTECTION_MODE         : integer := 31;
			FLASH_SEQ_READ_DATA_COUNT           : integer := 2;
			FLASH_ADDR_ALIGNMENT_BITS           : integer := 1;
			FLASH_READ_CYCLE_MAX_INDEX          : integer := 4;
			FLASH_RESET_CYCLE_MAX_INDEX         : integer := 29;
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  : integer := 112;
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX : integer := 40603248;
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX : integer := 35382;
			PARALLEL_MODE                       : boolean := true;
			READ_AND_WRITE_MODE                 : boolean := true;
			WRAPPING_BURST_MODE                 : boolean := false;
			IS_DUAL_BOOT                        : string  := "False";
			IS_ERAM_SKIP                        : string  := "False";
			IS_COMPRESSED_IMAGE                 : string  := "False"
		);
		port (
			clock                   : in  std_logic                     := 'X';             -- clk
			reset_n                 : in  std_logic                     := 'X';             -- reset_n
			avmm_data_addr          : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			avmm_data_read          : in  std_logic                     := 'X';             -- read
			avmm_data_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_data_write         : in  std_logic                     := 'X';             -- write
			avmm_data_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avmm_data_waitrequest   : out std_logic;                                        -- waitrequest
			avmm_data_readdatavalid : out std_logic;                                        -- readdatavalid
			avmm_data_burstcount    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			avmm_csr_addr           : in  std_logic                     := 'X';             -- address
			avmm_csr_read           : in  std_logic                     := 'X';             -- read
			avmm_csr_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_csr_write          : in  std_logic                     := 'X';             -- write
			avmm_csr_readdata       : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component altera_onchip_flash;

	component lms_ctr_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component lms_ctr_onchip_memory2_0;

	component lms_ctr_switch is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component lms_ctr_switch;

	component lms_ctr_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component lms_ctr_sysid_qsys_0;

	component lms_ctr_vctcxo_tamer_0_ctrl is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component lms_ctr_vctcxo_tamer_0_ctrl;

	component altera_customins_master_translator is
		generic (
			SHARED_COMB_AND_MULTI : integer := 0
		);
		port (
			ci_slave_dataa            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result           : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n                : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra           : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb           : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc          : in  std_logic                     := 'X';             -- writerc
			ci_slave_a                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c                : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus          : in  std_logic                     := 'X';             -- estatus
			comb_ci_master_dataa      : out std_logic_vector(31 downto 0);                    -- dataa
			comb_ci_master_datab      : out std_logic_vector(31 downto 0);                    -- datab
			comb_ci_master_result     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			comb_ci_master_n          : out std_logic_vector(7 downto 0);                     -- n
			comb_ci_master_readra     : out std_logic;                                        -- readra
			comb_ci_master_readrb     : out std_logic;                                        -- readrb
			comb_ci_master_writerc    : out std_logic;                                        -- writerc
			comb_ci_master_a          : out std_logic_vector(4 downto 0);                     -- a
			comb_ci_master_b          : out std_logic_vector(4 downto 0);                     -- b
			comb_ci_master_c          : out std_logic_vector(4 downto 0);                     -- c
			comb_ci_master_ipending   : out std_logic_vector(31 downto 0);                    -- ipending
			comb_ci_master_estatus    : out std_logic;                                        -- estatus
			ci_slave_multi_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_multi_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_multi_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_multi_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_multi_start      : in  std_logic                     := 'X';             -- start
			ci_slave_multi_done       : out std_logic;                                        -- done
			ci_slave_multi_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_dataa
			ci_slave_multi_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- multi_datab
			ci_slave_multi_result     : out std_logic_vector(31 downto 0);                    -- multi_result
			ci_slave_multi_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- multi_n
			ci_slave_multi_readra     : in  std_logic                     := 'X';             -- multi_readra
			ci_slave_multi_readrb     : in  std_logic                     := 'X';             -- multi_readrb
			ci_slave_multi_writerc    : in  std_logic                     := 'X';             -- multi_writerc
			ci_slave_multi_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_a
			ci_slave_multi_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_b
			ci_slave_multi_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- multi_c
			multi_ci_master_clk       : out std_logic;                                        -- clk
			multi_ci_master_reset     : out std_logic;                                        -- reset
			multi_ci_master_clken     : out std_logic;                                        -- clk_en
			multi_ci_master_reset_req : out std_logic;                                        -- reset_req
			multi_ci_master_start     : out std_logic;                                        -- start
			multi_ci_master_done      : in  std_logic                     := 'X';             -- done
			multi_ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			multi_ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			multi_ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			multi_ci_master_n         : out std_logic_vector(7 downto 0);                     -- n
			multi_ci_master_readra    : out std_logic;                                        -- readra
			multi_ci_master_readrb    : out std_logic;                                        -- readrb
			multi_ci_master_writerc   : out std_logic;                                        -- writerc
			multi_ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			multi_ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			multi_ci_master_c         : out std_logic_vector(4 downto 0)                      -- c
		);
	end component altera_customins_master_translator;

	component lms_ctr_nios2_cpu_custom_instruction_master_comb_xconnect is
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra     : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb     : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             -- writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             -- estatus
			ci_master0_dataa    : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master0_datab    : out std_logic_vector(31 downto 0);                    -- datab
			ci_master0_result   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master0_n        : out std_logic_vector(7 downto 0);                     -- n
			ci_master0_readra   : out std_logic;                                        -- readra
			ci_master0_readrb   : out std_logic;                                        -- readrb
			ci_master0_writerc  : out std_logic;                                        -- writerc
			ci_master0_a        : out std_logic_vector(4 downto 0);                     -- a
			ci_master0_b        : out std_logic_vector(4 downto 0);                     -- b
			ci_master0_c        : out std_logic_vector(4 downto 0);                     -- c
			ci_master0_ipending : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master0_estatus  : out std_logic                                         -- estatus
		);
	end component lms_ctr_nios2_cpu_custom_instruction_master_comb_xconnect;

	component altera_customins_slave_translator is
		generic (
			N_WIDTH          : integer := 8;
			USE_DONE         : integer := 1;
			NUM_FIXED_CYCLES : integer := 2
		);
		port (
			ci_slave_dataa      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- dataa
			ci_slave_datab      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- datab
			ci_slave_result     : out std_logic_vector(31 downto 0);                    -- result
			ci_slave_n          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- n
			ci_slave_readra     : in  std_logic                     := 'X';             -- readra
			ci_slave_readrb     : in  std_logic                     := 'X';             -- readrb
			ci_slave_writerc    : in  std_logic                     := 'X';             -- writerc
			ci_slave_a          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- a
			ci_slave_b          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- b
			ci_slave_c          : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- c
			ci_slave_ipending   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- ipending
			ci_slave_estatus    : in  std_logic                     := 'X';             -- estatus
			ci_master_dataa     : out std_logic_vector(31 downto 0);                    -- dataa
			ci_master_datab     : out std_logic_vector(31 downto 0);                    -- datab
			ci_master_result    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- result
			ci_master_n         : out std_logic_vector(7 downto 0);                     -- n
			ci_master_readra    : out std_logic;                                        -- readra
			ci_master_readrb    : out std_logic;                                        -- readrb
			ci_master_writerc   : out std_logic;                                        -- writerc
			ci_master_a         : out std_logic_vector(4 downto 0);                     -- a
			ci_master_b         : out std_logic_vector(4 downto 0);                     -- b
			ci_master_c         : out std_logic_vector(4 downto 0);                     -- c
			ci_master_ipending  : out std_logic_vector(31 downto 0);                    -- ipending
			ci_master_estatus   : out std_logic;                                        -- estatus
			ci_master_clk       : out std_logic;                                        -- clk
			ci_master_clken     : out std_logic;                                        -- clk_en
			ci_master_reset_req : out std_logic;                                        -- reset_req
			ci_master_reset     : out std_logic;                                        -- reset
			ci_master_start     : out std_logic;                                        -- start
			ci_master_done      : in  std_logic                     := 'X';             -- done
			ci_slave_clk        : in  std_logic                     := 'X';             -- clk
			ci_slave_clken      : in  std_logic                     := 'X';             -- clk_en
			ci_slave_reset_req  : in  std_logic                     := 'X';             -- reset_req
			ci_slave_reset      : in  std_logic                     := 'X';             -- reset
			ci_slave_start      : in  std_logic                     := 'X';             -- start
			ci_slave_done       : out std_logic                                         -- done
		);
	end component altera_customins_slave_translator;

	component lms_ctr_mm_interconnect_0 is
		port (
			clk_main_clk_clk                               : in  std_logic                     := 'X';             -- clk
			dual_boot_0_nreset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			nios2_cpu_reset_reset_bridge_in_reset_reset    : in  std_logic                     := 'X';             -- reset
			nios2_cpu_data_master_address                  : in  std_logic_vector(21 downto 0) := (others => 'X'); -- address
			nios2_cpu_data_master_waitrequest              : out std_logic;                                        -- waitrequest
			nios2_cpu_data_master_byteenable               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_cpu_data_master_read                     : in  std_logic                     := 'X';             -- read
			nios2_cpu_data_master_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_cpu_data_master_write                    : in  std_logic                     := 'X';             -- write
			nios2_cpu_data_master_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_cpu_data_master_debugaccess              : in  std_logic                     := 'X';             -- debugaccess
			nios2_cpu_instruction_master_address           : in  std_logic_vector(21 downto 0) := (others => 'X'); -- address
			nios2_cpu_instruction_master_waitrequest       : out std_logic;                                        -- waitrequest
			nios2_cpu_instruction_master_read              : in  std_logic                     := 'X';             -- read
			nios2_cpu_instruction_master_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			Av_FIFO_Int_0_avalon_slave_0_address           : out std_logic_vector(1 downto 0);                     -- address
			Av_FIFO_Int_0_avalon_slave_0_write             : out std_logic;                                        -- write
			Av_FIFO_Int_0_avalon_slave_0_read              : out std_logic;                                        -- read
			Av_FIFO_Int_0_avalon_slave_0_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Av_FIFO_Int_0_avalon_slave_0_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			Av_FIFO_Int_0_avalon_slave_0_chipselect        : out std_logic;                                        -- chipselect
			Avalon_MM_external_0_avs_s0_address            : out std_logic_vector(7 downto 0);                     -- address
			Avalon_MM_external_0_avs_s0_write              : out std_logic;                                        -- write
			Avalon_MM_external_0_avs_s0_read               : out std_logic;                                        -- read
			Avalon_MM_external_0_avs_s0_readdata           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			Avalon_MM_external_0_avs_s0_writedata          : out std_logic_vector(7 downto 0);                     -- writedata
			Avalon_MM_external_0_avs_s0_readdatavalid      : in  std_logic                     := 'X';             -- readdatavalid
			Avalon_MM_external_0_avs_s0_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			dac_spi_spi_control_port_address               : out std_logic_vector(2 downto 0);                     -- address
			dac_spi_spi_control_port_write                 : out std_logic;                                        -- write
			dac_spi_spi_control_port_read                  : out std_logic;                                        -- read
			dac_spi_spi_control_port_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			dac_spi_spi_control_port_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			dac_spi_spi_control_port_chipselect            : out std_logic;                                        -- chipselect
			dual_boot_0_avalon_address                     : out std_logic_vector(2 downto 0);                     -- address
			dual_boot_0_avalon_write                       : out std_logic;                                        -- write
			dual_boot_0_avalon_read                        : out std_logic;                                        -- read
			dual_boot_0_avalon_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dual_boot_0_avalon_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			flash_spi_spi_control_port_address             : out std_logic_vector(2 downto 0);                     -- address
			flash_spi_spi_control_port_write               : out std_logic;                                        -- write
			flash_spi_spi_control_port_read                : out std_logic;                                        -- read
			flash_spi_spi_control_port_readdata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			flash_spi_spi_control_port_writedata           : out std_logic_vector(15 downto 0);                    -- writedata
			flash_spi_spi_control_port_chipselect          : out std_logic;                                        -- chipselect
			fpga_spi_spi_control_port_address              : out std_logic_vector(2 downto 0);                     -- address
			fpga_spi_spi_control_port_write                : out std_logic;                                        -- write
			fpga_spi_spi_control_port_read                 : out std_logic;                                        -- read
			fpga_spi_spi_control_port_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			fpga_spi_spi_control_port_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			fpga_spi_spi_control_port_chipselect           : out std_logic;                                        -- chipselect
			i2c_opencores_0_avalon_slave_0_address         : out std_logic_vector(2 downto 0);                     -- address
			i2c_opencores_0_avalon_slave_0_write           : out std_logic;                                        -- write
			i2c_opencores_0_avalon_slave_0_readdata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			i2c_opencores_0_avalon_slave_0_writedata       : out std_logic_vector(7 downto 0);                     -- writedata
			i2c_opencores_0_avalon_slave_0_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			i2c_opencores_0_avalon_slave_0_chipselect      : out std_logic;                                        -- chipselect
			leds_s1_address                                : out std_logic_vector(1 downto 0);                     -- address
			leds_s1_write                                  : out std_logic;                                        -- write
			leds_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_s1_writedata                              : out std_logic_vector(31 downto 0);                    -- writedata
			leds_s1_chipselect                             : out std_logic;                                        -- chipselect
			lms_ctr_gpio_s1_address                        : out std_logic_vector(2 downto 0);                     -- address
			lms_ctr_gpio_s1_write                          : out std_logic;                                        -- write
			lms_ctr_gpio_s1_readdata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			lms_ctr_gpio_s1_writedata                      : out std_logic_vector(31 downto 0);                    -- writedata
			lms_ctr_gpio_s1_chipselect                     : out std_logic;                                        -- chipselect
			nios2_cpu_debug_mem_slave_address              : out std_logic_vector(8 downto 0);                     -- address
			nios2_cpu_debug_mem_slave_write                : out std_logic;                                        -- write
			nios2_cpu_debug_mem_slave_read                 : out std_logic;                                        -- read
			nios2_cpu_debug_mem_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_cpu_debug_mem_slave_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_cpu_debug_mem_slave_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_cpu_debug_mem_slave_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			nios2_cpu_debug_mem_slave_debugaccess          : out std_logic;                                        -- debugaccess
			onchip_flash_0_csr_address                     : out std_logic_vector(0 downto 0);                     -- address
			onchip_flash_0_csr_write                       : out std_logic;                                        -- write
			onchip_flash_0_csr_read                        : out std_logic;                                        -- read
			onchip_flash_0_csr_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_flash_0_csr_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_flash_0_data_address                    : out std_logic_vector(17 downto 0);                    -- address
			onchip_flash_0_data_write                      : out std_logic;                                        -- write
			onchip_flash_0_data_read                       : out std_logic;                                        -- read
			onchip_flash_0_data_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_flash_0_data_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_flash_0_data_burstcount                 : out std_logic_vector(3 downto 0);                     -- burstcount
			onchip_flash_0_data_readdatavalid              : in  std_logic                     := 'X';             -- readdatavalid
			onchip_flash_0_data_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			onchip_memory2_0_s1_address                    : out std_logic_vector(9 downto 0);                     -- address
			onchip_memory2_0_s1_write                      : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                 : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                      : out std_logic;                                        -- clken
			switch_s1_address                              : out std_logic_vector(1 downto 0);                     -- address
			switch_s1_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_qsys_0_control_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			vctcxo_tamer_0_ctrl_s1_address                 : out std_logic_vector(1 downto 0);                     -- address
			vctcxo_tamer_0_ctrl_s1_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component lms_ctr_mm_interconnect_0;

	component lms_ctr_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component lms_ctr_irq_mapper;

	component lms_ctr_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lms_ctr_rst_controller;

	component lms_ctr_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component lms_ctr_rst_controller_001;

	signal nios2_cpu_custom_instruction_master_readra                                  : std_logic;                     -- nios2_cpu:D_ci_readra -> nios2_cpu_custom_instruction_master_translator:ci_slave_readra
	signal nios2_cpu_custom_instruction_master_a                                       : std_logic_vector(4 downto 0);  -- nios2_cpu:D_ci_a -> nios2_cpu_custom_instruction_master_translator:ci_slave_a
	signal nios2_cpu_custom_instruction_master_b                                       : std_logic_vector(4 downto 0);  -- nios2_cpu:D_ci_b -> nios2_cpu_custom_instruction_master_translator:ci_slave_b
	signal nios2_cpu_custom_instruction_master_c                                       : std_logic_vector(4 downto 0);  -- nios2_cpu:D_ci_c -> nios2_cpu_custom_instruction_master_translator:ci_slave_c
	signal nios2_cpu_custom_instruction_master_readrb                                  : std_logic;                     -- nios2_cpu:D_ci_readrb -> nios2_cpu_custom_instruction_master_translator:ci_slave_readrb
	signal nios2_cpu_custom_instruction_master_ipending                                : std_logic_vector(31 downto 0); -- nios2_cpu:W_ci_ipending -> nios2_cpu_custom_instruction_master_translator:ci_slave_ipending
	signal nios2_cpu_custom_instruction_master_n                                       : std_logic_vector(7 downto 0);  -- nios2_cpu:D_ci_n -> nios2_cpu_custom_instruction_master_translator:ci_slave_n
	signal nios2_cpu_custom_instruction_master_result                                  : std_logic_vector(31 downto 0); -- nios2_cpu_custom_instruction_master_translator:ci_slave_result -> nios2_cpu:E_ci_result
	signal nios2_cpu_custom_instruction_master_estatus                                 : std_logic;                     -- nios2_cpu:W_ci_estatus -> nios2_cpu_custom_instruction_master_translator:ci_slave_estatus
	signal nios2_cpu_custom_instruction_master_datab                                   : std_logic_vector(31 downto 0); -- nios2_cpu:E_ci_datab -> nios2_cpu_custom_instruction_master_translator:ci_slave_datab
	signal nios2_cpu_custom_instruction_master_dataa                                   : std_logic_vector(31 downto 0); -- nios2_cpu:E_ci_dataa -> nios2_cpu_custom_instruction_master_translator:ci_slave_dataa
	signal nios2_cpu_custom_instruction_master_writerc                                 : std_logic;                     -- nios2_cpu:D_ci_writerc -> nios2_cpu_custom_instruction_master_translator:ci_slave_writerc
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_result        : std_logic_vector(31 downto 0); -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_cpu_custom_instruction_master_translator:comb_ci_master_result
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra        : std_logic;                     -- nios2_cpu_custom_instruction_master_translator:comb_ci_master_readra -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_readra
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_a             : std_logic_vector(4 downto 0);  -- nios2_cpu_custom_instruction_master_translator:comb_ci_master_a -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_a
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_b             : std_logic_vector(4 downto 0);  -- nios2_cpu_custom_instruction_master_translator:comb_ci_master_b -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_b
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb        : std_logic;                     -- nios2_cpu_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_readrb
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_c             : std_logic_vector(4 downto 0);  -- nios2_cpu_custom_instruction_master_translator:comb_ci_master_c -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_c
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus       : std_logic;                     -- nios2_cpu_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_estatus
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending      : std_logic_vector(31 downto 0); -- nios2_cpu_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_ipending
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab         : std_logic_vector(31 downto 0); -- nios2_cpu_custom_instruction_master_translator:comb_ci_master_datab -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_datab
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa         : std_logic_vector(31 downto 0); -- nios2_cpu_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_dataa
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc       : std_logic;                     -- nios2_cpu_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_writerc
	signal nios2_cpu_custom_instruction_master_translator_comb_ci_master_n             : std_logic_vector(7 downto 0);  -- nios2_cpu_custom_instruction_master_translator:comb_ci_master_n -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_slave_n
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result         : std_logic_vector(31 downto 0); -- nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_result
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra         : std_logic;                     -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a              : std_logic_vector(4 downto 0);  -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_a
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b              : std_logic_vector(4 downto 0);  -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_b
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb         : std_logic;                     -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c              : std_logic_vector(4 downto 0);  -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_c
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus        : std_logic;                     -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending       : std_logic_vector(31 downto 0); -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab          : std_logic_vector(31 downto 0); -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa          : std_logic_vector(31 downto 0); -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc        : std_logic;                     -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	signal nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n              : std_logic_vector(7 downto 0);  -- nios2_cpu_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_slave_n
	signal nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result : std_logic_vector(31 downto 0); -- nios_custom_instr_bitswap_0:result -> nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_result
	signal nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab  : std_logic_vector(31 downto 0); -- nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_datab -> nios_custom_instr_bitswap_0:datab
	signal nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa  : std_logic_vector(31 downto 0); -- nios2_cpu_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> nios_custom_instr_bitswap_0:dataa
	signal nios2_cpu_data_master_readdata                                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	signal nios2_cpu_data_master_waitrequest                                           : std_logic;                     -- mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	signal nios2_cpu_data_master_debugaccess                                           : std_logic;                     -- nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	signal nios2_cpu_data_master_address                                               : std_logic_vector(21 downto 0); -- nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	signal nios2_cpu_data_master_byteenable                                            : std_logic_vector(3 downto 0);  -- nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	signal nios2_cpu_data_master_read                                                  : std_logic;                     -- nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	signal nios2_cpu_data_master_write                                                 : std_logic;                     -- nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	signal nios2_cpu_data_master_writedata                                             : std_logic_vector(31 downto 0); -- nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	signal nios2_cpu_instruction_master_readdata                                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	signal nios2_cpu_instruction_master_waitrequest                                    : std_logic;                     -- mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	signal nios2_cpu_instruction_master_address                                        : std_logic_vector(21 downto 0); -- nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	signal nios2_cpu_instruction_master_read                                           : std_logic;                     -- nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	signal mm_interconnect_0_dual_boot_0_avalon_readdata                               : std_logic_vector(31 downto 0); -- dual_boot_0:avmm_rcv_readdata -> mm_interconnect_0:dual_boot_0_avalon_readdata
	signal mm_interconnect_0_dual_boot_0_avalon_address                                : std_logic_vector(2 downto 0);  -- mm_interconnect_0:dual_boot_0_avalon_address -> dual_boot_0:avmm_rcv_address
	signal mm_interconnect_0_dual_boot_0_avalon_read                                   : std_logic;                     -- mm_interconnect_0:dual_boot_0_avalon_read -> dual_boot_0:avmm_rcv_read
	signal mm_interconnect_0_dual_boot_0_avalon_write                                  : std_logic;                     -- mm_interconnect_0:dual_boot_0_avalon_write -> dual_boot_0:avmm_rcv_write
	signal mm_interconnect_0_dual_boot_0_avalon_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:dual_boot_0_avalon_writedata -> dual_boot_0:avmm_rcv_writedata
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect                   : std_logic;                     -- mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_chipselect -> Av_FIFO_Int_0:chipselect
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata                     : std_logic_vector(31 downto 0); -- Av_FIFO_Int_0:readdata -> mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_readdata
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_address -> Av_FIFO_Int_0:address
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read                         : std_logic;                     -- mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_read -> Av_FIFO_Int_0:read
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write                        : std_logic;                     -- mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_write -> Av_FIFO_Int_0:write
	signal mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_writedata -> Av_FIFO_Int_0:writedata
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect                 : std_logic;                     -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_chipselect -> i2c_opencores_0:wb_stb_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata                   : std_logic_vector(7 downto 0);  -- i2c_opencores_0:wb_dat_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_readdata
	signal i2c_opencores_0_avalon_slave_0_waitrequest                                  : std_logic;                     -- i2c_opencores_0:wb_ack_o -> i2c_opencores_0_avalon_slave_0_waitrequest:in
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address                    : std_logic_vector(2 downto 0);  -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_address -> i2c_opencores_0:wb_adr_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write                      : std_logic;                     -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_write -> i2c_opencores_0:wb_we_i
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata                  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:i2c_opencores_0_avalon_slave_0_writedata -> i2c_opencores_0:wb_dat_i
	signal mm_interconnect_0_avalon_mm_external_0_avs_s0_readdata                      : std_logic_vector(7 downto 0);  -- Avalon_MM_external_0:avs_s0_readdata -> mm_interconnect_0:Avalon_MM_external_0_avs_s0_readdata
	signal mm_interconnect_0_avalon_mm_external_0_avs_s0_waitrequest                   : std_logic;                     -- Avalon_MM_external_0:avs_s0_waitrequest -> mm_interconnect_0:Avalon_MM_external_0_avs_s0_waitrequest
	signal mm_interconnect_0_avalon_mm_external_0_avs_s0_address                       : std_logic_vector(7 downto 0);  -- mm_interconnect_0:Avalon_MM_external_0_avs_s0_address -> Avalon_MM_external_0:avs_s0_address
	signal mm_interconnect_0_avalon_mm_external_0_avs_s0_read                          : std_logic;                     -- mm_interconnect_0:Avalon_MM_external_0_avs_s0_read -> Avalon_MM_external_0:avs_s0_read
	signal mm_interconnect_0_avalon_mm_external_0_avs_s0_readdatavalid                 : std_logic;                     -- Avalon_MM_external_0:avs_s0_readdatavalid -> mm_interconnect_0:Avalon_MM_external_0_avs_s0_readdatavalid
	signal mm_interconnect_0_avalon_mm_external_0_avs_s0_write                         : std_logic;                     -- mm_interconnect_0:Avalon_MM_external_0_avs_s0_write -> Avalon_MM_external_0:avs_s0_write
	signal mm_interconnect_0_avalon_mm_external_0_avs_s0_writedata                     : std_logic_vector(7 downto 0);  -- mm_interconnect_0:Avalon_MM_external_0_avs_s0_writedata -> Avalon_MM_external_0:avs_s0_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata                       : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                        : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_onchip_flash_0_csr_readdata                               : std_logic_vector(31 downto 0); -- onchip_flash_0:avmm_csr_readdata -> mm_interconnect_0:onchip_flash_0_csr_readdata
	signal mm_interconnect_0_onchip_flash_0_csr_address                                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:onchip_flash_0_csr_address -> onchip_flash_0:avmm_csr_addr
	signal mm_interconnect_0_onchip_flash_0_csr_read                                   : std_logic;                     -- mm_interconnect_0:onchip_flash_0_csr_read -> onchip_flash_0:avmm_csr_read
	signal mm_interconnect_0_onchip_flash_0_csr_write                                  : std_logic;                     -- mm_interconnect_0:onchip_flash_0_csr_write -> onchip_flash_0:avmm_csr_write
	signal mm_interconnect_0_onchip_flash_0_csr_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_flash_0_csr_writedata -> onchip_flash_0:avmm_csr_writedata
	signal mm_interconnect_0_onchip_flash_0_data_readdata                              : std_logic_vector(31 downto 0); -- onchip_flash_0:avmm_data_readdata -> mm_interconnect_0:onchip_flash_0_data_readdata
	signal mm_interconnect_0_onchip_flash_0_data_waitrequest                           : std_logic;                     -- onchip_flash_0:avmm_data_waitrequest -> mm_interconnect_0:onchip_flash_0_data_waitrequest
	signal mm_interconnect_0_onchip_flash_0_data_address                               : std_logic_vector(17 downto 0); -- mm_interconnect_0:onchip_flash_0_data_address -> onchip_flash_0:avmm_data_addr
	signal mm_interconnect_0_onchip_flash_0_data_read                                  : std_logic;                     -- mm_interconnect_0:onchip_flash_0_data_read -> onchip_flash_0:avmm_data_read
	signal mm_interconnect_0_onchip_flash_0_data_readdatavalid                         : std_logic;                     -- onchip_flash_0:avmm_data_readdatavalid -> mm_interconnect_0:onchip_flash_0_data_readdatavalid
	signal mm_interconnect_0_onchip_flash_0_data_write                                 : std_logic;                     -- mm_interconnect_0:onchip_flash_0_data_write -> onchip_flash_0:avmm_data_write
	signal mm_interconnect_0_onchip_flash_0_data_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_flash_0_data_writedata -> onchip_flash_0:avmm_data_writedata
	signal mm_interconnect_0_onchip_flash_0_data_burstcount                            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_flash_0_data_burstcount -> onchip_flash_0:avmm_data_burstcount
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata                        : std_logic_vector(31 downto 0); -- nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest                     : std_logic;                     -- nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess                     : std_logic;                     -- mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_address                         : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_read                            : std_logic;                     -- mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_write                           : std_logic;                     -- mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	signal mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_switch_s1_readdata                                        : std_logic_vector(31 downto 0); -- switch:readdata -> mm_interconnect_0:switch_s1_readdata
	signal mm_interconnect_0_switch_s1_address                                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_s1_address -> switch:address
	signal mm_interconnect_0_leds_s1_chipselect                                        : std_logic;                     -- mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	signal mm_interconnect_0_leds_s1_readdata                                          : std_logic_vector(31 downto 0); -- leds:readdata -> mm_interconnect_0:leds_s1_readdata
	signal mm_interconnect_0_leds_s1_address                                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_s1_address -> leds:address
	signal mm_interconnect_0_leds_s1_write                                             : std_logic;                     -- mm_interconnect_0:leds_s1_write -> mm_interconnect_0_leds_s1_write:in
	signal mm_interconnect_0_leds_s1_writedata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_s1_writedata -> leds:writedata
	signal mm_interconnect_0_lms_ctr_gpio_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:lms_ctr_gpio_s1_chipselect -> lms_ctr_gpio:chipselect
	signal mm_interconnect_0_lms_ctr_gpio_s1_readdata                                  : std_logic_vector(31 downto 0); -- lms_ctr_gpio:readdata -> mm_interconnect_0:lms_ctr_gpio_s1_readdata
	signal mm_interconnect_0_lms_ctr_gpio_s1_address                                   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:lms_ctr_gpio_s1_address -> lms_ctr_gpio:address
	signal mm_interconnect_0_lms_ctr_gpio_s1_write                                     : std_logic;                     -- mm_interconnect_0:lms_ctr_gpio_s1_write -> mm_interconnect_0_lms_ctr_gpio_s1_write:in
	signal mm_interconnect_0_lms_ctr_gpio_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:lms_ctr_gpio_s1_writedata -> lms_ctr_gpio:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                              : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                               : std_logic_vector(9 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                                 : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                                 : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_vctcxo_tamer_0_ctrl_s1_readdata                           : std_logic_vector(31 downto 0); -- vctcxo_tamer_0_ctrl:readdata -> mm_interconnect_0:vctcxo_tamer_0_ctrl_s1_readdata
	signal mm_interconnect_0_vctcxo_tamer_0_ctrl_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:vctcxo_tamer_0_ctrl_s1_address -> vctcxo_tamer_0_ctrl:address
	signal mm_interconnect_0_fpga_spi_spi_control_port_chipselect                      : std_logic;                     -- mm_interconnect_0:fpga_spi_spi_control_port_chipselect -> fpga_spi:spi_select
	signal mm_interconnect_0_fpga_spi_spi_control_port_readdata                        : std_logic_vector(15 downto 0); -- fpga_spi:data_to_cpu -> mm_interconnect_0:fpga_spi_spi_control_port_readdata
	signal mm_interconnect_0_fpga_spi_spi_control_port_address                         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:fpga_spi_spi_control_port_address -> fpga_spi:mem_addr
	signal mm_interconnect_0_fpga_spi_spi_control_port_read                            : std_logic;                     -- mm_interconnect_0:fpga_spi_spi_control_port_read -> mm_interconnect_0_fpga_spi_spi_control_port_read:in
	signal mm_interconnect_0_fpga_spi_spi_control_port_write                           : std_logic;                     -- mm_interconnect_0:fpga_spi_spi_control_port_write -> mm_interconnect_0_fpga_spi_spi_control_port_write:in
	signal mm_interconnect_0_fpga_spi_spi_control_port_writedata                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:fpga_spi_spi_control_port_writedata -> fpga_spi:data_from_cpu
	signal mm_interconnect_0_dac_spi_spi_control_port_chipselect                       : std_logic;                     -- mm_interconnect_0:dac_spi_spi_control_port_chipselect -> dac_spi:spi_select
	signal mm_interconnect_0_dac_spi_spi_control_port_readdata                         : std_logic_vector(15 downto 0); -- dac_spi:data_to_cpu -> mm_interconnect_0:dac_spi_spi_control_port_readdata
	signal mm_interconnect_0_dac_spi_spi_control_port_address                          : std_logic_vector(2 downto 0);  -- mm_interconnect_0:dac_spi_spi_control_port_address -> dac_spi:mem_addr
	signal mm_interconnect_0_dac_spi_spi_control_port_read                             : std_logic;                     -- mm_interconnect_0:dac_spi_spi_control_port_read -> mm_interconnect_0_dac_spi_spi_control_port_read:in
	signal mm_interconnect_0_dac_spi_spi_control_port_write                            : std_logic;                     -- mm_interconnect_0:dac_spi_spi_control_port_write -> mm_interconnect_0_dac_spi_spi_control_port_write:in
	signal mm_interconnect_0_dac_spi_spi_control_port_writedata                        : std_logic_vector(15 downto 0); -- mm_interconnect_0:dac_spi_spi_control_port_writedata -> dac_spi:data_from_cpu
	signal mm_interconnect_0_flash_spi_spi_control_port_chipselect                     : std_logic;                     -- mm_interconnect_0:flash_spi_spi_control_port_chipselect -> flash_spi:spi_select
	signal mm_interconnect_0_flash_spi_spi_control_port_readdata                       : std_logic_vector(15 downto 0); -- flash_spi:data_to_cpu -> mm_interconnect_0:flash_spi_spi_control_port_readdata
	signal mm_interconnect_0_flash_spi_spi_control_port_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:flash_spi_spi_control_port_address -> flash_spi:mem_addr
	signal mm_interconnect_0_flash_spi_spi_control_port_read                           : std_logic;                     -- mm_interconnect_0:flash_spi_spi_control_port_read -> mm_interconnect_0_flash_spi_spi_control_port_read:in
	signal mm_interconnect_0_flash_spi_spi_control_port_write                          : std_logic;                     -- mm_interconnect_0:flash_spi_spi_control_port_write -> mm_interconnect_0_flash_spi_spi_control_port_write:in
	signal mm_interconnect_0_flash_spi_spi_control_port_writedata                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:flash_spi_spi_control_port_writedata -> flash_spi:data_from_cpu
	signal irq_mapper_receiver0_irq                                                    : std_logic;                     -- i2c_opencores_0:wb_inta_o -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                    : std_logic;                     -- fpga_spi:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                    : std_logic;                     -- dac_spi:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                    : std_logic;                     -- flash_spi:irq -> irq_mapper:receiver3_irq
	signal nios2_cpu_irq_irq                                                           : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_cpu:irq
	signal rst_controller_reset_out_reset                                              : std_logic;                     -- rst_controller:reset_out -> [Avalon_MM_external_0:reset_reset, i2c_opencores_0:wb_rst_i, irq_mapper:reset, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                          : std_logic;                     -- rst_controller:reset_req -> [nios2_cpu:reset_req, rst_translator:reset_req_in]
	signal nios2_cpu_debug_reset_request_reset                                         : std_logic;                     -- nios2_cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in0]
	signal rst_controller_001_reset_out_reset                                          : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:dual_boot_0_nreset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_001_reset_out_reset:in, rst_translator_001:in_reset]
	signal rst_controller_001_reset_out_reset_req                                      : std_logic;                     -- rst_controller_001:reset_req -> [onchip_memory2_0:reset_req, rst_translator_001:reset_req_in]
	signal reset_reset_n_ports_inv                                                     : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv                        : std_logic;                     -- i2c_opencores_0_avalon_slave_0_waitrequest:inv -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_waitrequest
	signal mm_interconnect_0_leds_s1_write_ports_inv                                   : std_logic;                     -- mm_interconnect_0_leds_s1_write:inv -> leds:write_n
	signal mm_interconnect_0_lms_ctr_gpio_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_lms_ctr_gpio_s1_write:inv -> lms_ctr_gpio:write_n
	signal mm_interconnect_0_fpga_spi_spi_control_port_read_ports_inv                  : std_logic;                     -- mm_interconnect_0_fpga_spi_spi_control_port_read:inv -> fpga_spi:read_n
	signal mm_interconnect_0_fpga_spi_spi_control_port_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_fpga_spi_spi_control_port_write:inv -> fpga_spi:write_n
	signal mm_interconnect_0_dac_spi_spi_control_port_read_ports_inv                   : std_logic;                     -- mm_interconnect_0_dac_spi_spi_control_port_read:inv -> dac_spi:read_n
	signal mm_interconnect_0_dac_spi_spi_control_port_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_dac_spi_spi_control_port_write:inv -> dac_spi:write_n
	signal mm_interconnect_0_flash_spi_spi_control_port_read_ports_inv                 : std_logic;                     -- mm_interconnect_0_flash_spi_spi_control_port_read:inv -> flash_spi:read_n
	signal mm_interconnect_0_flash_spi_spi_control_port_write_ports_inv                : std_logic;                     -- mm_interconnect_0_flash_spi_spi_control_port_write:inv -> flash_spi:write_n
	signal rst_controller_reset_out_reset_ports_inv                                    : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Av_FIFO_Int_0:rsi_nrst, dac_spi:reset_n, flash_spi:reset_n, fpga_spi:reset_n, leds:reset_n, lms_ctr_gpio:reset_n, nios2_cpu:reset_n, switch:reset_n, sysid_qsys_0:reset_n, vctcxo_tamer_0_ctrl:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                                : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [dual_boot_0:nreset, onchip_flash_0:reset_n]

begin

	av_fifo_int_0 : component avfifo
		generic map (
			width => 32
		)
		port map (
			clk            => clk_clk,                                                   --          clock.clk
			address        => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address,    -- avalon_slave_0.address
			chipselect     => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect, --               .chipselect
			write          => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write,      --               .write
			writedata      => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata,  --               .writedata
			read           => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read,       --               .read
			readdata       => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata,   --               .readdata
			rsi_nrst       => rst_controller_reset_out_reset_ports_inv,                  --          reset.reset_n
			coe_if_d       => exfifo_if_d_export,                                        --       cnd_if_d.export
			coe_if_rd      => exfifo_if_rd_export,                                       --      cnd_if_rd.export
			coe_of_wrfull  => exfifo_of_wrfull_export,                                   --  cnd_of_wrfull.export
			coe_of_wr      => exfifo_of_wr_export,                                       --      cnd_of_wr.export
			coe_of_d       => exfifo_of_d_export,                                        --       cnd_of_d.export
			coe_if_rdempty => exfifo_if_rdempty_export,                                  -- cnd_if_rdempty.export
			coe_fifo_rst   => exfifo_rst_export                                          --   cnd_fifo_rst.export
		);

	avalon_mm_external_0 : component Avalon_MM_external
		port map (
			avs_s0_address       => mm_interconnect_0_avalon_mm_external_0_avs_s0_address,       --       avs_s0.address
			avs_s0_read          => mm_interconnect_0_avalon_mm_external_0_avs_s0_read,          --             .read
			avs_s0_readdata      => mm_interconnect_0_avalon_mm_external_0_avs_s0_readdata,      --             .readdata
			avs_s0_write         => mm_interconnect_0_avalon_mm_external_0_avs_s0_write,         --             .write
			avs_s0_writedata     => mm_interconnect_0_avalon_mm_external_0_avs_s0_writedata,     --             .writedata
			avs_s0_waitrequest   => mm_interconnect_0_avalon_mm_external_0_avs_s0_waitrequest,   --             .waitrequest
			avs_s0_readdatavalid => mm_interconnect_0_avalon_mm_external_0_avs_s0_readdatavalid, --             .readdatavalid
			clock_clk            => clk_clk,                                                     --        clock.clk
			reset_reset          => rst_controller_reset_out_reset,                              --        reset.reset
			avm_m0_address       => avm_m0_address,                                              --       avm_m0.address
			avm_m0_read          => avm_m0_read,                                                 --             .read
			avm_m0_waitrequest   => avm_m0_waitrequest,                                          --             .waitrequest
			avm_m0_readdata      => avm_m0_readdata,                                             --             .readdata
			avm_m0_write         => avm_m0_write,                                                --             .write
			avm_m0_writedata     => avm_m0_writedata,                                            --             .writedata
			avm_m0_readdatavalid => avm_m0_readdatavalid,                                        --             .readdatavalid
			clock_source_clk     => avm_m0_clk_clk,                                              -- clock_source.clk
			reset_source_reset   => avm_m0_reset_reset                                           -- reset_source.reset
		);

	dac_spi : component lms_ctr_dac_spi
		port map (
			clk           => clk_clk,                                                    --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                   --            reset.reset_n
			data_from_cpu => mm_interconnect_0_dac_spi_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_dac_spi_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_dac_spi_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_dac_spi_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_dac_spi_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_dac_spi_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver2_irq,                                   --              irq.irq
			MISO          => dac_spi_ext_MISO,                                           --         external.export
			MOSI          => dac_spi_ext_MOSI,                                           --                 .export
			SCLK          => dac_spi_ext_SCLK,                                           --                 .export
			SS_n          => dac_spi_ext_SS_n                                            --                 .export
		);

	dual_boot_0 : component altera_dual_boot
		generic map (
			INTENDED_DEVICE_FAMILY => "MAX 10",
			CONFIG_CYCLE           => 15,
			RESET_TIMER_CYCLE      => 21
		)
		port map (
			clk                => clk_clk,                                        --    clk.clk
			nreset             => rst_controller_001_reset_out_reset_ports_inv,   -- nreset.reset_n
			avmm_rcv_address   => mm_interconnect_0_dual_boot_0_avalon_address,   -- avalon.address
			avmm_rcv_read      => mm_interconnect_0_dual_boot_0_avalon_read,      --       .read
			avmm_rcv_writedata => mm_interconnect_0_dual_boot_0_avalon_writedata, --       .writedata
			avmm_rcv_write     => mm_interconnect_0_dual_boot_0_avalon_write,     --       .write
			avmm_rcv_readdata  => mm_interconnect_0_dual_boot_0_avalon_readdata   --       .readdata
		);

	flash_spi : component lms_ctr_flash_spi
		port map (
			clk           => clk_clk,                                                      --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                     --            reset.reset_n
			data_from_cpu => mm_interconnect_0_flash_spi_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_flash_spi_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_flash_spi_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_flash_spi_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_flash_spi_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_flash_spi_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver3_irq,                                     --              irq.irq
			MISO          => flash_spi_MISO,                                               --         external.export
			MOSI          => flash_spi_MOSI,                                               --                 .export
			SCLK          => flash_spi_SCLK,                                               --                 .export
			SS_n          => flash_spi_SS_n                                                --                 .export
		);

	fpga_spi : component lms_ctr_fpga_spi
		port map (
			clk           => clk_clk,                                                     --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                    --            reset.reset_n
			data_from_cpu => mm_interconnect_0_fpga_spi_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_fpga_spi_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_fpga_spi_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_fpga_spi_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_fpga_spi_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_fpga_spi_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver1_irq,                                    --              irq.irq
			MISO          => fpga_spi_ext_MISO,                                           --         external.export
			MOSI          => fpga_spi_ext_MOSI,                                           --                 .export
			SCLK          => fpga_spi_ext_SCLK,                                           --                 .export
			SS_n          => fpga_spi_ext_SS_n                                            --                 .export
		);

	i2c_opencores_0 : component i2c_opencores
		port map (
			wb_clk_i   => clk_clk,                                                     --            clock.clk
			wb_rst_i   => rst_controller_reset_out_reset,                              --      clock_reset.reset
			scl_pad_io => i2c_scl_export,                                              --       export_scl.export
			sda_pad_io => i2c_sda_export,                                              --       export_sda.export
			wb_adr_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address,    --   avalon_slave_0.address
			wb_dat_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata,  --                 .writedata
			wb_dat_o   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata,   --                 .readdata
			wb_we_i    => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write,      --                 .write
			wb_stb_i   => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect, --                 .chipselect
			wb_ack_o   => i2c_opencores_0_avalon_slave_0_waitrequest,                  --                 .waitrequest_n
			wb_inta_o  => irq_mapper_receiver0_irq                                     -- interrupt_sender.irq
		);

	leds : component lms_ctr_leds
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_s1_readdata,        --                    .readdata
			out_port   => leds_external_connection_export            -- external_connection.export
		);

	lms_ctr_gpio : component lms_ctr_lms_ctr_gpio
		port map (
			clk        => clk_clk,                                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_lms_ctr_gpio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_lms_ctr_gpio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_lms_ctr_gpio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_lms_ctr_gpio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_lms_ctr_gpio_s1_readdata,        --                    .readdata
			out_port   => lms_ctr_gpio_external_connection_export            -- external_connection.export
		);

	nios2_cpu : component lms_ctr_nios2_cpu
		port map (
			clk                                 => clk_clk,                                                 --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                      --                          .reset_req
			d_address                           => nios2_cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_cpu_data_master_read,                              --                          .read
			d_readdata                          => nios2_cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_cpu_data_master_write,                             --                          .write
			d_writedata                         => nios2_cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_cpu_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata,   --                          .writedata
			E_ci_result                         => nios2_cpu_custom_instruction_master_result,              -- custom_instruction_master.result
			D_ci_a                              => nios2_cpu_custom_instruction_master_a,                   --                          .a
			D_ci_b                              => nios2_cpu_custom_instruction_master_b,                   --                          .b
			D_ci_c                              => nios2_cpu_custom_instruction_master_c,                   --                          .c
			D_ci_n                              => nios2_cpu_custom_instruction_master_n,                   --                          .n
			D_ci_readra                         => nios2_cpu_custom_instruction_master_readra,              --                          .readra
			D_ci_readrb                         => nios2_cpu_custom_instruction_master_readrb,              --                          .readrb
			D_ci_writerc                        => nios2_cpu_custom_instruction_master_writerc,             --                          .writerc
			E_ci_dataa                          => nios2_cpu_custom_instruction_master_dataa,               --                          .dataa
			E_ci_datab                          => nios2_cpu_custom_instruction_master_datab,               --                          .datab
			E_ci_multi_clock                    => open,                                                    --                          .clk
			E_ci_multi_reset                    => open,                                                    --                          .reset
			E_ci_multi_reset_req                => open,                                                    --                          .reset_req
			W_ci_estatus                        => nios2_cpu_custom_instruction_master_estatus,             --                          .estatus
			W_ci_ipending                       => nios2_cpu_custom_instruction_master_ipending             --                          .ipending
		);

	nios_custom_instr_bitswap_0 : component bitswap_qsys
		port map (
			dataa  => nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa,  -- s1.dataa
			datab  => nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab,  --   .datab
			result => nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result  --   .result
		);

	onchip_flash_0 : component altera_onchip_flash
		generic map (
			INIT_FILENAME                       => "lms_ctr_onchip_flash_0.hex",
			INIT_FILENAME_SIM                   => "lms_ctr_onchip_flash_0.dat",
			DEVICE_FAMILY                       => "MAX 10",
			PART_NAME                           => "10M16SAU169C8G",
			DEVICE_ID                           => "16",
			SECTOR1_START_ADDR                  => 0,
			SECTOR1_END_ADDR                    => 4095,
			SECTOR2_START_ADDR                  => 4096,
			SECTOR2_END_ADDR                    => 8191,
			SECTOR3_START_ADDR                  => 8192,
			SECTOR3_END_ADDR                    => 47103,
			SECTOR4_START_ADDR                  => 47104,
			SECTOR4_END_ADDR                    => 75775,
			SECTOR5_START_ADDR                  => 75776,
			SECTOR5_END_ADDR                    => 143359,
			MIN_VALID_ADDR                      => 0,
			MAX_VALID_ADDR                      => 143359,
			MIN_UFM_VALID_ADDR                  => 0,
			MAX_UFM_VALID_ADDR                  => 8191,
			SECTOR1_MAP                         => 1,
			SECTOR2_MAP                         => 2,
			SECTOR3_MAP                         => 3,
			SECTOR4_MAP                         => 4,
			SECTOR5_MAP                         => 5,
			ADDR_RANGE1_END_ADDR                => 143359,
			ADDR_RANGE2_END_ADDR                => 143359,
			ADDR_RANGE1_OFFSET                  => 1024,
			ADDR_RANGE2_OFFSET                  => 0,
			ADDR_RANGE3_OFFSET                  => 0,
			AVMM_DATA_ADDR_WIDTH                => 18,
			AVMM_DATA_DATA_WIDTH                => 32,
			AVMM_DATA_BURSTCOUNT_WIDTH          => 4,
			SECTOR_READ_PROTECTION_MODE         => 1,
			FLASH_SEQ_READ_DATA_COUNT           => 4,
			FLASH_ADDR_ALIGNMENT_BITS           => 2,
			FLASH_READ_CYCLE_MAX_INDEX          => 4,
			FLASH_RESET_CYCLE_MAX_INDEX         => 7,
			FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  => 36,
			FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX => 10752027,
			FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX => 9369,
			PARALLEL_MODE                       => true,
			READ_AND_WRITE_MODE                 => true,
			WRAPPING_BURST_MODE                 => false,
			IS_DUAL_BOOT                        => "True",
			IS_ERAM_SKIP                        => "True",
			IS_COMPRESSED_IMAGE                 => "True"
		)
		port map (
			clock                   => clk_clk,                                             --    clk.clk
			reset_n                 => rst_controller_001_reset_out_reset_ports_inv,        -- nreset.reset_n
			avmm_data_addr          => mm_interconnect_0_onchip_flash_0_data_address,       --   data.address
			avmm_data_read          => mm_interconnect_0_onchip_flash_0_data_read,          --       .read
			avmm_data_writedata     => mm_interconnect_0_onchip_flash_0_data_writedata,     --       .writedata
			avmm_data_write         => mm_interconnect_0_onchip_flash_0_data_write,         --       .write
			avmm_data_readdata      => mm_interconnect_0_onchip_flash_0_data_readdata,      --       .readdata
			avmm_data_waitrequest   => mm_interconnect_0_onchip_flash_0_data_waitrequest,   --       .waitrequest
			avmm_data_readdatavalid => mm_interconnect_0_onchip_flash_0_data_readdatavalid, --       .readdatavalid
			avmm_data_burstcount    => mm_interconnect_0_onchip_flash_0_data_burstcount,    --       .burstcount
			avmm_csr_addr           => mm_interconnect_0_onchip_flash_0_csr_address(0),     --    csr.address
			avmm_csr_read           => mm_interconnect_0_onchip_flash_0_csr_read,           --       .read
			avmm_csr_writedata      => mm_interconnect_0_onchip_flash_0_csr_writedata,      --       .writedata
			avmm_csr_write          => mm_interconnect_0_onchip_flash_0_csr_write,          --       .write
			avmm_csr_readdata       => mm_interconnect_0_onchip_flash_0_csr_readdata        --       .readdata
		);

	onchip_memory2_0 : component lms_ctr_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,               -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,           --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	switch : component lms_ctr_switch
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switch_s1_address,      --                  s1.address
			readdata => mm_interconnect_0_switch_s1_readdata,     --                    .readdata
			in_port  => switch_external_connection_export         -- external_connection.export
		);

	sysid_qsys_0 : component lms_ctr_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	vctcxo_tamer_0_ctrl : component lms_ctr_vctcxo_tamer_0_ctrl
		port map (
			clk      => clk_clk,                                           --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address  => mm_interconnect_0_vctcxo_tamer_0_ctrl_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_vctcxo_tamer_0_ctrl_s1_readdata, --                    .readdata
			in_port  => vctcxo_tamer_0_ctrl_export                         -- external_connection.export
		);

	nios2_cpu_custom_instruction_master_translator : component altera_customins_master_translator
		generic map (
			SHARED_COMB_AND_MULTI => 1
		)
		port map (
			ci_slave_dataa            => nios2_cpu_custom_instruction_master_dataa,                              --       ci_slave.dataa
			ci_slave_datab            => nios2_cpu_custom_instruction_master_datab,                              --               .datab
			ci_slave_result           => nios2_cpu_custom_instruction_master_result,                             --               .result
			ci_slave_n                => nios2_cpu_custom_instruction_master_n,                                  --               .n
			ci_slave_readra           => nios2_cpu_custom_instruction_master_readra,                             --               .readra
			ci_slave_readrb           => nios2_cpu_custom_instruction_master_readrb,                             --               .readrb
			ci_slave_writerc          => nios2_cpu_custom_instruction_master_writerc,                            --               .writerc
			ci_slave_a                => nios2_cpu_custom_instruction_master_a,                                  --               .a
			ci_slave_b                => nios2_cpu_custom_instruction_master_b,                                  --               .b
			ci_slave_c                => nios2_cpu_custom_instruction_master_c,                                  --               .c
			ci_slave_ipending         => nios2_cpu_custom_instruction_master_ipending,                           --               .ipending
			ci_slave_estatus          => nios2_cpu_custom_instruction_master_estatus,                            --               .estatus
			comb_ci_master_dataa      => nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa,    -- comb_ci_master.dataa
			comb_ci_master_datab      => nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab,    --               .datab
			comb_ci_master_result     => nios2_cpu_custom_instruction_master_translator_comb_ci_master_result,   --               .result
			comb_ci_master_n          => nios2_cpu_custom_instruction_master_translator_comb_ci_master_n,        --               .n
			comb_ci_master_readra     => nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra,   --               .readra
			comb_ci_master_readrb     => nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb,   --               .readrb
			comb_ci_master_writerc    => nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc,  --               .writerc
			comb_ci_master_a          => nios2_cpu_custom_instruction_master_translator_comb_ci_master_a,        --               .a
			comb_ci_master_b          => nios2_cpu_custom_instruction_master_translator_comb_ci_master_b,        --               .b
			comb_ci_master_c          => nios2_cpu_custom_instruction_master_translator_comb_ci_master_c,        --               .c
			comb_ci_master_ipending   => nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending, --               .ipending
			comb_ci_master_estatus    => nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus,  --               .estatus
			ci_slave_multi_clk        => '0',                                                                    --    (terminated)
			ci_slave_multi_reset      => '0',                                                                    --    (terminated)
			ci_slave_multi_clken      => '0',                                                                    --    (terminated)
			ci_slave_multi_reset_req  => '0',                                                                    --    (terminated)
			ci_slave_multi_start      => '0',                                                                    --    (terminated)
			ci_slave_multi_done       => open,                                                                   --    (terminated)
			ci_slave_multi_dataa      => "00000000000000000000000000000000",                                     --    (terminated)
			ci_slave_multi_datab      => "00000000000000000000000000000000",                                     --    (terminated)
			ci_slave_multi_result     => open,                                                                   --    (terminated)
			ci_slave_multi_n          => "00000000",                                                             --    (terminated)
			ci_slave_multi_readra     => '0',                                                                    --    (terminated)
			ci_slave_multi_readrb     => '0',                                                                    --    (terminated)
			ci_slave_multi_writerc    => '0',                                                                    --    (terminated)
			ci_slave_multi_a          => "00000",                                                                --    (terminated)
			ci_slave_multi_b          => "00000",                                                                --    (terminated)
			ci_slave_multi_c          => "00000",                                                                --    (terminated)
			multi_ci_master_clk       => open,                                                                   --    (terminated)
			multi_ci_master_reset     => open,                                                                   --    (terminated)
			multi_ci_master_clken     => open,                                                                   --    (terminated)
			multi_ci_master_reset_req => open,                                                                   --    (terminated)
			multi_ci_master_start     => open,                                                                   --    (terminated)
			multi_ci_master_done      => '0',                                                                    --    (terminated)
			multi_ci_master_dataa     => open,                                                                   --    (terminated)
			multi_ci_master_datab     => open,                                                                   --    (terminated)
			multi_ci_master_result    => "00000000000000000000000000000000",                                     --    (terminated)
			multi_ci_master_n         => open,                                                                   --    (terminated)
			multi_ci_master_readra    => open,                                                                   --    (terminated)
			multi_ci_master_readrb    => open,                                                                   --    (terminated)
			multi_ci_master_writerc   => open,                                                                   --    (terminated)
			multi_ci_master_a         => open,                                                                   --    (terminated)
			multi_ci_master_b         => open,                                                                   --    (terminated)
			multi_ci_master_c         => open                                                                    --    (terminated)
		);

	nios2_cpu_custom_instruction_master_comb_xconnect : component lms_ctr_nios2_cpu_custom_instruction_master_comb_xconnect
		port map (
			ci_slave_dataa      => nios2_cpu_custom_instruction_master_translator_comb_ci_master_dataa,    --   ci_slave.dataa
			ci_slave_datab      => nios2_cpu_custom_instruction_master_translator_comb_ci_master_datab,    --           .datab
			ci_slave_result     => nios2_cpu_custom_instruction_master_translator_comb_ci_master_result,   --           .result
			ci_slave_n          => nios2_cpu_custom_instruction_master_translator_comb_ci_master_n,        --           .n
			ci_slave_readra     => nios2_cpu_custom_instruction_master_translator_comb_ci_master_readra,   --           .readra
			ci_slave_readrb     => nios2_cpu_custom_instruction_master_translator_comb_ci_master_readrb,   --           .readrb
			ci_slave_writerc    => nios2_cpu_custom_instruction_master_translator_comb_ci_master_writerc,  --           .writerc
			ci_slave_a          => nios2_cpu_custom_instruction_master_translator_comb_ci_master_a,        --           .a
			ci_slave_b          => nios2_cpu_custom_instruction_master_translator_comb_ci_master_b,        --           .b
			ci_slave_c          => nios2_cpu_custom_instruction_master_translator_comb_ci_master_c,        --           .c
			ci_slave_ipending   => nios2_cpu_custom_instruction_master_translator_comb_ci_master_ipending, --           .ipending
			ci_slave_estatus    => nios2_cpu_custom_instruction_master_translator_comb_ci_master_estatus,  --           .estatus
			ci_master0_dataa    => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa,     -- ci_master0.dataa
			ci_master0_datab    => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab,     --           .datab
			ci_master0_result   => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result,    --           .result
			ci_master0_n        => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n,         --           .n
			ci_master0_readra   => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra,    --           .readra
			ci_master0_readrb   => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb,    --           .readrb
			ci_master0_writerc  => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc,   --           .writerc
			ci_master0_a        => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a,         --           .a
			ci_master0_b        => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b,         --           .b
			ci_master0_c        => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c,         --           .c
			ci_master0_ipending => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending,  --           .ipending
			ci_master0_estatus  => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus    --           .estatus
		);

	nios2_cpu_custom_instruction_master_comb_slave_translator0 : component altera_customins_slave_translator
		generic map (
			N_WIDTH          => 8,
			USE_DONE         => 0,
			NUM_FIXED_CYCLES => 1
		)
		port map (
			ci_slave_dataa      => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_dataa,          --  ci_slave.dataa
			ci_slave_datab      => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_datab,          --          .datab
			ci_slave_result     => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_result,         --          .result
			ci_slave_n          => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_n,              --          .n
			ci_slave_readra     => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readra,         --          .readra
			ci_slave_readrb     => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_readrb,         --          .readrb
			ci_slave_writerc    => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_writerc,        --          .writerc
			ci_slave_a          => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_a,              --          .a
			ci_slave_b          => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_b,              --          .b
			ci_slave_c          => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_c,              --          .c
			ci_slave_ipending   => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_ipending,       --          .ipending
			ci_slave_estatus    => nios2_cpu_custom_instruction_master_comb_xconnect_ci_master0_estatus,        --          .estatus
			ci_master_dataa     => nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_dataa,  -- ci_master.dataa
			ci_master_datab     => nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_datab,  --          .datab
			ci_master_result    => nios2_cpu_custom_instruction_master_comb_slave_translator0_ci_master_result, --          .result
			ci_master_n         => open,                                                                        -- (terminated)
			ci_master_readra    => open,                                                                        -- (terminated)
			ci_master_readrb    => open,                                                                        -- (terminated)
			ci_master_writerc   => open,                                                                        -- (terminated)
			ci_master_a         => open,                                                                        -- (terminated)
			ci_master_b         => open,                                                                        -- (terminated)
			ci_master_c         => open,                                                                        -- (terminated)
			ci_master_ipending  => open,                                                                        -- (terminated)
			ci_master_estatus   => open,                                                                        -- (terminated)
			ci_master_clk       => open,                                                                        -- (terminated)
			ci_master_clken     => open,                                                                        -- (terminated)
			ci_master_reset_req => open,                                                                        -- (terminated)
			ci_master_reset     => open,                                                                        -- (terminated)
			ci_master_start     => open,                                                                        -- (terminated)
			ci_master_done      => '0',                                                                         -- (terminated)
			ci_slave_clk        => '0',                                                                         -- (terminated)
			ci_slave_clken      => '0',                                                                         -- (terminated)
			ci_slave_reset_req  => '0',                                                                         -- (terminated)
			ci_slave_reset      => '0',                                                                         -- (terminated)
			ci_slave_start      => '0',                                                                         -- (terminated)
			ci_slave_done       => open                                                                         -- (terminated)
		);

	mm_interconnect_0 : component lms_ctr_mm_interconnect_0
		port map (
			clk_main_clk_clk                               => clk_clk,                                                     --                             clk_main_clk.clk
			dual_boot_0_nreset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                          -- dual_boot_0_nreset_reset_bridge_in_reset.reset
			nios2_cpu_reset_reset_bridge_in_reset_reset    => rst_controller_reset_out_reset,                              --    nios2_cpu_reset_reset_bridge_in_reset.reset
			nios2_cpu_data_master_address                  => nios2_cpu_data_master_address,                               --                    nios2_cpu_data_master.address
			nios2_cpu_data_master_waitrequest              => nios2_cpu_data_master_waitrequest,                           --                                         .waitrequest
			nios2_cpu_data_master_byteenable               => nios2_cpu_data_master_byteenable,                            --                                         .byteenable
			nios2_cpu_data_master_read                     => nios2_cpu_data_master_read,                                  --                                         .read
			nios2_cpu_data_master_readdata                 => nios2_cpu_data_master_readdata,                              --                                         .readdata
			nios2_cpu_data_master_write                    => nios2_cpu_data_master_write,                                 --                                         .write
			nios2_cpu_data_master_writedata                => nios2_cpu_data_master_writedata,                             --                                         .writedata
			nios2_cpu_data_master_debugaccess              => nios2_cpu_data_master_debugaccess,                           --                                         .debugaccess
			nios2_cpu_instruction_master_address           => nios2_cpu_instruction_master_address,                        --             nios2_cpu_instruction_master.address
			nios2_cpu_instruction_master_waitrequest       => nios2_cpu_instruction_master_waitrequest,                    --                                         .waitrequest
			nios2_cpu_instruction_master_read              => nios2_cpu_instruction_master_read,                           --                                         .read
			nios2_cpu_instruction_master_readdata          => nios2_cpu_instruction_master_readdata,                       --                                         .readdata
			Av_FIFO_Int_0_avalon_slave_0_address           => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address,      --             Av_FIFO_Int_0_avalon_slave_0.address
			Av_FIFO_Int_0_avalon_slave_0_write             => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write,        --                                         .write
			Av_FIFO_Int_0_avalon_slave_0_read              => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read,         --                                         .read
			Av_FIFO_Int_0_avalon_slave_0_readdata          => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata,     --                                         .readdata
			Av_FIFO_Int_0_avalon_slave_0_writedata         => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata,    --                                         .writedata
			Av_FIFO_Int_0_avalon_slave_0_chipselect        => mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect,   --                                         .chipselect
			Avalon_MM_external_0_avs_s0_address            => mm_interconnect_0_avalon_mm_external_0_avs_s0_address,       --              Avalon_MM_external_0_avs_s0.address
			Avalon_MM_external_0_avs_s0_write              => mm_interconnect_0_avalon_mm_external_0_avs_s0_write,         --                                         .write
			Avalon_MM_external_0_avs_s0_read               => mm_interconnect_0_avalon_mm_external_0_avs_s0_read,          --                                         .read
			Avalon_MM_external_0_avs_s0_readdata           => mm_interconnect_0_avalon_mm_external_0_avs_s0_readdata,      --                                         .readdata
			Avalon_MM_external_0_avs_s0_writedata          => mm_interconnect_0_avalon_mm_external_0_avs_s0_writedata,     --                                         .writedata
			Avalon_MM_external_0_avs_s0_readdatavalid      => mm_interconnect_0_avalon_mm_external_0_avs_s0_readdatavalid, --                                         .readdatavalid
			Avalon_MM_external_0_avs_s0_waitrequest        => mm_interconnect_0_avalon_mm_external_0_avs_s0_waitrequest,   --                                         .waitrequest
			dac_spi_spi_control_port_address               => mm_interconnect_0_dac_spi_spi_control_port_address,          --                 dac_spi_spi_control_port.address
			dac_spi_spi_control_port_write                 => mm_interconnect_0_dac_spi_spi_control_port_write,            --                                         .write
			dac_spi_spi_control_port_read                  => mm_interconnect_0_dac_spi_spi_control_port_read,             --                                         .read
			dac_spi_spi_control_port_readdata              => mm_interconnect_0_dac_spi_spi_control_port_readdata,         --                                         .readdata
			dac_spi_spi_control_port_writedata             => mm_interconnect_0_dac_spi_spi_control_port_writedata,        --                                         .writedata
			dac_spi_spi_control_port_chipselect            => mm_interconnect_0_dac_spi_spi_control_port_chipselect,       --                                         .chipselect
			dual_boot_0_avalon_address                     => mm_interconnect_0_dual_boot_0_avalon_address,                --                       dual_boot_0_avalon.address
			dual_boot_0_avalon_write                       => mm_interconnect_0_dual_boot_0_avalon_write,                  --                                         .write
			dual_boot_0_avalon_read                        => mm_interconnect_0_dual_boot_0_avalon_read,                   --                                         .read
			dual_boot_0_avalon_readdata                    => mm_interconnect_0_dual_boot_0_avalon_readdata,               --                                         .readdata
			dual_boot_0_avalon_writedata                   => mm_interconnect_0_dual_boot_0_avalon_writedata,              --                                         .writedata
			flash_spi_spi_control_port_address             => mm_interconnect_0_flash_spi_spi_control_port_address,        --               flash_spi_spi_control_port.address
			flash_spi_spi_control_port_write               => mm_interconnect_0_flash_spi_spi_control_port_write,          --                                         .write
			flash_spi_spi_control_port_read                => mm_interconnect_0_flash_spi_spi_control_port_read,           --                                         .read
			flash_spi_spi_control_port_readdata            => mm_interconnect_0_flash_spi_spi_control_port_readdata,       --                                         .readdata
			flash_spi_spi_control_port_writedata           => mm_interconnect_0_flash_spi_spi_control_port_writedata,      --                                         .writedata
			flash_spi_spi_control_port_chipselect          => mm_interconnect_0_flash_spi_spi_control_port_chipselect,     --                                         .chipselect
			fpga_spi_spi_control_port_address              => mm_interconnect_0_fpga_spi_spi_control_port_address,         --                fpga_spi_spi_control_port.address
			fpga_spi_spi_control_port_write                => mm_interconnect_0_fpga_spi_spi_control_port_write,           --                                         .write
			fpga_spi_spi_control_port_read                 => mm_interconnect_0_fpga_spi_spi_control_port_read,            --                                         .read
			fpga_spi_spi_control_port_readdata             => mm_interconnect_0_fpga_spi_spi_control_port_readdata,        --                                         .readdata
			fpga_spi_spi_control_port_writedata            => mm_interconnect_0_fpga_spi_spi_control_port_writedata,       --                                         .writedata
			fpga_spi_spi_control_port_chipselect           => mm_interconnect_0_fpga_spi_spi_control_port_chipselect,      --                                         .chipselect
			i2c_opencores_0_avalon_slave_0_address         => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address,    --           i2c_opencores_0_avalon_slave_0.address
			i2c_opencores_0_avalon_slave_0_write           => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write,      --                                         .write
			i2c_opencores_0_avalon_slave_0_readdata        => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata,   --                                         .readdata
			i2c_opencores_0_avalon_slave_0_writedata       => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata,  --                                         .writedata
			i2c_opencores_0_avalon_slave_0_waitrequest     => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv,        --                                         .waitrequest
			i2c_opencores_0_avalon_slave_0_chipselect      => mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect, --                                         .chipselect
			leds_s1_address                                => mm_interconnect_0_leds_s1_address,                           --                                  leds_s1.address
			leds_s1_write                                  => mm_interconnect_0_leds_s1_write,                             --                                         .write
			leds_s1_readdata                               => mm_interconnect_0_leds_s1_readdata,                          --                                         .readdata
			leds_s1_writedata                              => mm_interconnect_0_leds_s1_writedata,                         --                                         .writedata
			leds_s1_chipselect                             => mm_interconnect_0_leds_s1_chipselect,                        --                                         .chipselect
			lms_ctr_gpio_s1_address                        => mm_interconnect_0_lms_ctr_gpio_s1_address,                   --                          lms_ctr_gpio_s1.address
			lms_ctr_gpio_s1_write                          => mm_interconnect_0_lms_ctr_gpio_s1_write,                     --                                         .write
			lms_ctr_gpio_s1_readdata                       => mm_interconnect_0_lms_ctr_gpio_s1_readdata,                  --                                         .readdata
			lms_ctr_gpio_s1_writedata                      => mm_interconnect_0_lms_ctr_gpio_s1_writedata,                 --                                         .writedata
			lms_ctr_gpio_s1_chipselect                     => mm_interconnect_0_lms_ctr_gpio_s1_chipselect,                --                                         .chipselect
			nios2_cpu_debug_mem_slave_address              => mm_interconnect_0_nios2_cpu_debug_mem_slave_address,         --                nios2_cpu_debug_mem_slave.address
			nios2_cpu_debug_mem_slave_write                => mm_interconnect_0_nios2_cpu_debug_mem_slave_write,           --                                         .write
			nios2_cpu_debug_mem_slave_read                 => mm_interconnect_0_nios2_cpu_debug_mem_slave_read,            --                                         .read
			nios2_cpu_debug_mem_slave_readdata             => mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata,        --                                         .readdata
			nios2_cpu_debug_mem_slave_writedata            => mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata,       --                                         .writedata
			nios2_cpu_debug_mem_slave_byteenable           => mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable,      --                                         .byteenable
			nios2_cpu_debug_mem_slave_waitrequest          => mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest,     --                                         .waitrequest
			nios2_cpu_debug_mem_slave_debugaccess          => mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess,     --                                         .debugaccess
			onchip_flash_0_csr_address                     => mm_interconnect_0_onchip_flash_0_csr_address,                --                       onchip_flash_0_csr.address
			onchip_flash_0_csr_write                       => mm_interconnect_0_onchip_flash_0_csr_write,                  --                                         .write
			onchip_flash_0_csr_read                        => mm_interconnect_0_onchip_flash_0_csr_read,                   --                                         .read
			onchip_flash_0_csr_readdata                    => mm_interconnect_0_onchip_flash_0_csr_readdata,               --                                         .readdata
			onchip_flash_0_csr_writedata                   => mm_interconnect_0_onchip_flash_0_csr_writedata,              --                                         .writedata
			onchip_flash_0_data_address                    => mm_interconnect_0_onchip_flash_0_data_address,               --                      onchip_flash_0_data.address
			onchip_flash_0_data_write                      => mm_interconnect_0_onchip_flash_0_data_write,                 --                                         .write
			onchip_flash_0_data_read                       => mm_interconnect_0_onchip_flash_0_data_read,                  --                                         .read
			onchip_flash_0_data_readdata                   => mm_interconnect_0_onchip_flash_0_data_readdata,              --                                         .readdata
			onchip_flash_0_data_writedata                  => mm_interconnect_0_onchip_flash_0_data_writedata,             --                                         .writedata
			onchip_flash_0_data_burstcount                 => mm_interconnect_0_onchip_flash_0_data_burstcount,            --                                         .burstcount
			onchip_flash_0_data_readdatavalid              => mm_interconnect_0_onchip_flash_0_data_readdatavalid,         --                                         .readdatavalid
			onchip_flash_0_data_waitrequest                => mm_interconnect_0_onchip_flash_0_data_waitrequest,           --                                         .waitrequest
			onchip_memory2_0_s1_address                    => mm_interconnect_0_onchip_memory2_0_s1_address,               --                      onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                      => mm_interconnect_0_onchip_memory2_0_s1_write,                 --                                         .write
			onchip_memory2_0_s1_readdata                   => mm_interconnect_0_onchip_memory2_0_s1_readdata,              --                                         .readdata
			onchip_memory2_0_s1_writedata                  => mm_interconnect_0_onchip_memory2_0_s1_writedata,             --                                         .writedata
			onchip_memory2_0_s1_byteenable                 => mm_interconnect_0_onchip_memory2_0_s1_byteenable,            --                                         .byteenable
			onchip_memory2_0_s1_chipselect                 => mm_interconnect_0_onchip_memory2_0_s1_chipselect,            --                                         .chipselect
			onchip_memory2_0_s1_clken                      => mm_interconnect_0_onchip_memory2_0_s1_clken,                 --                                         .clken
			switch_s1_address                              => mm_interconnect_0_switch_s1_address,                         --                                switch_s1.address
			switch_s1_readdata                             => mm_interconnect_0_switch_s1_readdata,                        --                                         .readdata
			sysid_qsys_0_control_slave_address             => mm_interconnect_0_sysid_qsys_0_control_slave_address,        --               sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata            => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,       --                                         .readdata
			vctcxo_tamer_0_ctrl_s1_address                 => mm_interconnect_0_vctcxo_tamer_0_ctrl_s1_address,            --                   vctcxo_tamer_0_ctrl_s1.address
			vctcxo_tamer_0_ctrl_s1_readdata                => mm_interconnect_0_vctcxo_tamer_0_ctrl_s1_readdata            --                                         .readdata
		);

	irq_mapper : component lms_ctr_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => nios2_cpu_irq_irq               --    sender.irq
		);

	rst_controller : component lms_ctr_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,             -- reset_in0.reset
			reset_in1      => nios2_cpu_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,      -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,  --          .reset_req
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_in2      => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	rst_controller_001 : component lms_ctr_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => nios2_cpu_debug_reset_request_reset,    -- reset_in0.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_i2c_opencores_0_avalon_slave_0_inv <= not i2c_opencores_0_avalon_slave_0_waitrequest;

	mm_interconnect_0_leds_s1_write_ports_inv <= not mm_interconnect_0_leds_s1_write;

	mm_interconnect_0_lms_ctr_gpio_s1_write_ports_inv <= not mm_interconnect_0_lms_ctr_gpio_s1_write;

	mm_interconnect_0_fpga_spi_spi_control_port_read_ports_inv <= not mm_interconnect_0_fpga_spi_spi_control_port_read;

	mm_interconnect_0_fpga_spi_spi_control_port_write_ports_inv <= not mm_interconnect_0_fpga_spi_spi_control_port_write;

	mm_interconnect_0_dac_spi_spi_control_port_read_ports_inv <= not mm_interconnect_0_dac_spi_spi_control_port_read;

	mm_interconnect_0_dac_spi_spi_control_port_write_ports_inv <= not mm_interconnect_0_dac_spi_spi_control_port_write;

	mm_interconnect_0_flash_spi_spi_control_port_read_ports_inv <= not mm_interconnect_0_flash_spi_spi_control_port_read;

	mm_interconnect_0_flash_spi_spi_control_port_write_ports_inv <= not mm_interconnect_0_flash_spi_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of lms_ctr
